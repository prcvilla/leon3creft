leon3mp_original.vhd