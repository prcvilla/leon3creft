----------------------------------------------------------------------------
--  This file is a part of the GRLIB VHDL IP LIBRARY
--  Copyright (C) 2004 GAISLER RESEARCH
--
--  This program is free software; you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation; either version 2 of the License, or
--  (at your option) any later version.
--
--  See the file COPYING for the full details of the license.
--
-----------------------------------------------------------------------------
-- Entity: 	ahbrom
-- File:	ahbrom.vhd
-- Author:	Jiri Gaisler - Gaisler Research
-- Description:	AHB rom. 0/1-waitstate read
------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library grlib;
use grlib.amba.all;
use grlib.stdlib.all;
use grlib.devices.all;

entity ahbrom is
  generic (
    hindex  : integer := 0;
    haddr   : integer := 0;
    hmask   : integer := 16#fff#;
    pipe    : integer := 0;
    tech    : integer := 0;
    kbytes  : integer := 1);
  port (
    rst     : in  std_ulogic;
    clk     : in  std_ulogic;
    ahbsi   : in  ahb_slv_in_type;
    ahbso   : out ahb_slv_out_type
  );
end;

architecture rtl of ahbrom is
constant abits : integer := 9;
constant bytes : integer := 432;

constant hconfig : ahb_config_type := (
  0 => ahb_device_reg ( VENDOR_GAISLER, GAISLER_AHBROM, 0, 0, 0),
  4 => ahb_membar(haddr, '1', '1', hmask), others => zero32);

signal romdata : std_logic_vector(31 downto 0);
signal addr : std_logic_vector(abits-1 downto 2);
signal hsel, hready : std_ulogic;

begin

  ahbso.hresp   <= "00"; 
  ahbso.hsplit  <= (others => '0'); 
  ahbso.hirq    <= (others => '0');
  ahbso.hconfig <= hconfig;
  ahbso.hindex  <= hindex;

  reg : process (clk)
  begin
    if rising_edge(clk) then 
      addr <= ahbsi.haddr(abits-1 downto 2);
    end if;
  end process;

  p0 : if pipe = 0 generate
    ahbso.hrdata  <= ahbdrivedata(romdata);
    ahbso.hready  <= '1';
  end generate;

  p1 : if pipe = 1 generate
    reg2 : process (clk)
    begin
      if rising_edge(clk) then
	hsel <= ahbsi.hsel(hindex) and ahbsi.htrans(1);
	hready <= ahbsi.hready;
	ahbso.hready <=  (not rst) or (hsel and hready) or
	  (ahbsi.hsel(hindex) and not ahbsi.htrans(1) and ahbsi.hready);
	ahbso.hrdata  <= ahbdrivedata(romdata);
      end if;
    end process;
  end generate;

  comb : process (addr)
  begin
    case conv_integer(addr) is
	when 16#00000# => romdata <= X"0D100004";
when 16#00001# => romdata <= X"81C1A39C";
when 16#00002# => romdata <= X"01000000";
when 16#00003# => romdata <= X"9DE3BFC0";
when 16#00004# => romdata <= X"0510000A";
when 16#00005# => romdata <= X"8410A380";
when 16#00006# => romdata <= X"0710000B";
when 16#00007# => romdata <= X"8610E2F8";
when 16#00008# => romdata <= X"82100000";
when 16#00009# => romdata <= X"8620C002";
when 16#0000A# => romdata <= X"86A0E008";
when 16#0000B# => romdata <= X"36BFFFFF";
when 16#0000C# => romdata <= X"C0388003";
when 16#0000D# => romdata <= X"1110000B";
when 16#0000E# => romdata <= X"901222F8";
when 16#0000F# => romdata <= X"C0220000";
when 16#00010# => romdata <= X"400004CE";
when 16#00011# => romdata <= X"01000000";
when 16#00012# => romdata <= X"400004CE";
when 16#00013# => romdata <= X"01000000";
when 16#00014# => romdata <= X"4000050D";
when 16#00015# => romdata <= X"01000000";
when 16#00016# => romdata <= X"11100008";
when 16#00017# => romdata <= X"901223EC";
when 16#00018# => romdata <= X"40000481";
when 16#00019# => romdata <= X"01000000";
when 16#0001A# => romdata <= X"400008DA";
when 16#0001B# => romdata <= X"01000000";
when 16#0001C# => romdata <= X"400003A9";
when 16#0001D# => romdata <= X"01000000";
when 16#0001E# => romdata <= X"400004C4";
when 16#0001F# => romdata <= X"01000000";
when 16#00020# => romdata <= X"81C7E008";
when 16#00021# => romdata <= X"81E80000";
when 16#00022# => romdata <= X"9DE3BFA0";
when 16#00023# => romdata <= X"3B10000A";
when 16#00024# => romdata <= X"C20F6380";
when 16#00025# => romdata <= X"80A06000";
when 16#00026# => romdata <= X"12800022";
when 16#00027# => romdata <= X"3910000A";
when 16#00028# => romdata <= X"C2072384";
when 16#00029# => romdata <= X"35100008";
when 16#0002A# => romdata <= X"37100008";
when 16#0002B# => romdata <= X"B416A264";
when 16#0002C# => romdata <= X"B616E268";
when 16#0002D# => romdata <= X"B626C01A";
when 16#0002E# => romdata <= X"B73EE002";
when 16#0002F# => romdata <= X"B606FFFF";
when 16#00030# => romdata <= X"80A0401B";
when 16#00031# => romdata <= X"3A80000E";
when 16#00032# => romdata <= X"03000000";
when 16#00033# => romdata <= X"B8172384";
when 16#00034# => romdata <= X"82006001";
when 16#00035# => romdata <= X"85286002";
when 16#00036# => romdata <= X"C2270000";
when 16#00037# => romdata <= X"C2068002";
when 16#00038# => romdata <= X"9FC04000";
when 16#00039# => romdata <= X"01000000";
when 16#0003A# => romdata <= X"C2070000";
when 16#0003B# => romdata <= X"80A0401B";
when 16#0003C# => romdata <= X"0ABFFFF9";
when 16#0003D# => romdata <= X"82006001";
when 16#0003E# => romdata <= X"03000000";
when 16#0003F# => romdata <= X"82106000";
when 16#00040# => romdata <= X"80A06000";
when 16#00041# => romdata <= X"02800006";
when 16#00042# => romdata <= X"82102001";
when 16#00043# => romdata <= X"11100008";
when 16#00044# => romdata <= X"6FFFFFBC";
when 16#00045# => romdata <= X"90122240";
when 16#00046# => romdata <= X"82102001";
when 16#00047# => romdata <= X"C22F6380";
when 16#00048# => romdata <= X"81C7E008";
when 16#00049# => romdata <= X"81E80000";
when 16#0004A# => romdata <= X"9DE3BFA0";
when 16#0004B# => romdata <= X"81C7E008";
when 16#0004C# => romdata <= X"81E80000";
when 16#0004D# => romdata <= X"9DE3BFA0";
when 16#0004E# => romdata <= X"03000000";
when 16#0004F# => romdata <= X"82106000";
when 16#00050# => romdata <= X"80A06000";
when 16#00051# => romdata <= X"22800008";
when 16#00052# => romdata <= X"1110000B";
when 16#00053# => romdata <= X"11100008";
when 16#00054# => romdata <= X"1310000A";
when 16#00055# => romdata <= X"90122240";
when 16#00056# => romdata <= X"6FFFFFAA";
when 16#00057# => romdata <= X"92126388";
when 16#00058# => romdata <= X"1110000B";
when 16#00059# => romdata <= X"C20222F8";
when 16#0005A# => romdata <= X"80A06000";
when 16#0005B# => romdata <= X"02800009";
when 16#0005C# => romdata <= X"901222F8";
when 16#0005D# => romdata <= X"03000000";
when 16#0005E# => romdata <= X"82106000";
when 16#0005F# => romdata <= X"80A06000";
when 16#00060# => romdata <= X"02800004";
when 16#00061# => romdata <= X"01000000";
when 16#00062# => romdata <= X"9FC04000";
when 16#00063# => romdata <= X"01000000";
when 16#00064# => romdata <= X"81C7E008";
when 16#00065# => romdata <= X"81E80000";
when 16#00066# => romdata <= X"9DE3BFA0";
when 16#00067# => romdata <= X"81C7E008";
when 16#00068# => romdata <= X"81E80000";
when 16#00069# => romdata <= X"81C3E008";
when 16#0006A# => romdata <= X"01000000";
when 16#0006B# => romdata <= X"98120009";
when 16#0006C# => romdata <= X"81800008";
when 16#0006D# => romdata <= X"98880000";
when 16#0006E# => romdata <= X"99230009";
when 16#0006F# => romdata <= X"99230009";
when 16#00070# => romdata <= X"99230009";
when 16#00071# => romdata <= X"99230009";
when 16#00072# => romdata <= X"99230009";
when 16#00073# => romdata <= X"99230009";
when 16#00074# => romdata <= X"99230009";
when 16#00075# => romdata <= X"99230009";
when 16#00076# => romdata <= X"99230009";
when 16#00077# => romdata <= X"99230009";
when 16#00078# => romdata <= X"99230009";
when 16#00079# => romdata <= X"99230009";
when 16#0007A# => romdata <= X"99230009";
when 16#0007B# => romdata <= X"99230009";
when 16#0007C# => romdata <= X"99230009";
when 16#0007D# => romdata <= X"99230009";
when 16#0007E# => romdata <= X"99230009";
when 16#0007F# => romdata <= X"99230009";
when 16#00080# => romdata <= X"99230009";
when 16#00081# => romdata <= X"99230009";
when 16#00082# => romdata <= X"99230009";
when 16#00083# => romdata <= X"99230009";
when 16#00084# => romdata <= X"99230009";
when 16#00085# => romdata <= X"99230009";
when 16#00086# => romdata <= X"99230009";
when 16#00087# => romdata <= X"99230009";
when 16#00088# => romdata <= X"99230009";
when 16#00089# => romdata <= X"99230009";
when 16#0008A# => romdata <= X"99230009";
when 16#0008B# => romdata <= X"99230009";
when 16#0008C# => romdata <= X"99230009";
when 16#0008D# => romdata <= X"99230009";
when 16#0008E# => romdata <= X"99230000";
when 16#0008F# => romdata <= X"953A601F";
when 16#00090# => romdata <= X"940A000A";
when 16#00091# => romdata <= X"93400000";
when 16#00092# => romdata <= X"81C3E008";
when 16#00093# => romdata <= X"9083000A";
when 16#00094# => romdata <= X"9DE3BF98";
when 16#00095# => romdata <= X"F027A044";
when 16#00096# => romdata <= X"F227A048";
when 16#00097# => romdata <= X"F427A04C";
when 16#00098# => romdata <= X"C207A044";
when 16#00099# => romdata <= X"C4004000";
when 16#0009A# => romdata <= X"031FFFFF";
when 16#0009B# => romdata <= X"821063FF";
when 16#0009C# => romdata <= X"84088001";
when 16#0009D# => romdata <= X"C207A048";
when 16#0009E# => romdata <= X"C6004000";
when 16#0009F# => romdata <= X"031FFFFF";
when 16#000A0# => romdata <= X"821063FF";
when 16#000A1# => romdata <= X"8208C001";
when 16#000A2# => romdata <= X"90100002";
when 16#000A3# => romdata <= X"92100001";
when 16#000A4# => romdata <= X"7FFFFFC7";
when 16#000A5# => romdata <= X"01000000";
when 16#000A6# => romdata <= X"D03FBFF8";
when 16#000A7# => romdata <= X"C207BFF8";
when 16#000A8# => romdata <= X"83286010";
when 16#000A9# => romdata <= X"C407BFFC";
when 16#000AA# => romdata <= X"8530A010";
when 16#000AB# => romdata <= X"82108001";
when 16#000AC# => romdata <= X"C227BFFC";
when 16#000AD# => romdata <= X"C207BFF8";
when 16#000AE# => romdata <= X"83306010";
when 16#000AF# => romdata <= X"C227BFF8";
when 16#000B0# => romdata <= X"C407BFFC";
when 16#000B1# => romdata <= X"031FFFFF";
when 16#000B2# => romdata <= X"821063FF";
when 16#000B3# => romdata <= X"84088001";
when 16#000B4# => romdata <= X"C207A04C";
when 16#000B5# => romdata <= X"C4204000";
when 16#000B6# => romdata <= X"C207A044";
when 16#000B7# => romdata <= X"C2004000";
when 16#000B8# => romdata <= X"8330601F";
when 16#000B9# => romdata <= X"84100001";
when 16#000BA# => romdata <= X"C207A048";
when 16#000BB# => romdata <= X"C2004000";
when 16#000BC# => romdata <= X"8330601F";
when 16#000BD# => romdata <= X"82188001";
when 16#000BE# => romdata <= X"82086001";
when 16#000BF# => romdata <= X"84100001";
when 16#000C0# => romdata <= X"C207A04C";
when 16#000C1# => romdata <= X"8408A0FF";
when 16#000C2# => romdata <= X"8528A01F";
when 16#000C3# => romdata <= X"C8004000";
when 16#000C4# => romdata <= X"071FFFFF";
when 16#000C5# => romdata <= X"8610E3FF";
when 16#000C6# => romdata <= X"86090003";
when 16#000C7# => romdata <= X"8410C002";
when 16#000C8# => romdata <= X"C4204000";
when 16#000C9# => romdata <= X"81E80000";
when 16#000CA# => romdata <= X"81C3E008";
when 16#000CB# => romdata <= X"01000000";
when 16#000CC# => romdata <= X"9DE3BF60";
when 16#000CD# => romdata <= X"F027A044";
when 16#000CE# => romdata <= X"F227A048";
when 16#000CF# => romdata <= X"F427A04C";
when 16#000D0# => romdata <= X"C207A044";
when 16#000D1# => romdata <= X"C2004000";
when 16#000D2# => romdata <= X"B4102000";
when 16#000D3# => romdata <= X"B6100001";
when 16#000D4# => romdata <= X"B8102000";
when 16#000D5# => romdata <= X"3B1FFFFF";
when 16#000D6# => romdata <= X"BA1763FF";
when 16#000D7# => romdata <= X"B80E801C";
when 16#000D8# => romdata <= X"BA0EC01D";
when 16#000D9# => romdata <= X"F83FBFE0";
when 16#000DA# => romdata <= X"F81FBFE0";
when 16#000DB# => romdata <= X"BAA0001D";
when 16#000DC# => romdata <= X"B860001C";
when 16#000DD# => romdata <= X"F83FBFE8";
when 16#000DE# => romdata <= X"C207A048";
when 16#000DF# => romdata <= X"C2004000";
when 16#000E0# => romdata <= X"B4102000";
when 16#000E1# => romdata <= X"B6100001";
when 16#000E2# => romdata <= X"B8102000";
when 16#000E3# => romdata <= X"3B1FFFFF";
when 16#000E4# => romdata <= X"BA1763FF";
when 16#000E5# => romdata <= X"B80E801C";
when 16#000E6# => romdata <= X"BA0EC01D";
when 16#000E7# => romdata <= X"F83FBFD0";
when 16#000E8# => romdata <= X"F81FBFD0";
when 16#000E9# => romdata <= X"BAA0001D";
when 16#000EA# => romdata <= X"B860001C";
when 16#000EB# => romdata <= X"F83FBFD8";
when 16#000EC# => romdata <= X"C207A044";
when 16#000ED# => romdata <= X"C2004000";
when 16#000EE# => romdata <= X"8330601F";
when 16#000EF# => romdata <= X"820860FF";
when 16#000F0# => romdata <= X"83286003";
when 16#000F1# => romdata <= X"82078001";
when 16#000F2# => romdata <= X"F4187FE0";
when 16#000F3# => romdata <= X"C207A048";
when 16#000F4# => romdata <= X"C2004000";
when 16#000F5# => romdata <= X"8330601F";
when 16#000F6# => romdata <= X"820860FF";
when 16#000F7# => romdata <= X"83286003";
when 16#000F8# => romdata <= X"82078001";
when 16#000F9# => romdata <= X"F8187FD0";
when 16#000FA# => romdata <= X"BA86C01D";
when 16#000FB# => romdata <= X"B846801C";
when 16#000FC# => romdata <= X"F83FBFF8";
when 16#000FD# => romdata <= X"F81FBFF8";
when 16#000FE# => romdata <= X"8737201F";
when 16#000FF# => romdata <= X"84102000";
when 16#00100# => romdata <= X"C627BFF4";
when 16#00101# => romdata <= X"C41FBFF8";
when 16#00102# => romdata <= X"C43FBFC0";
when 16#00103# => romdata <= X"C41FBFF8";
when 16#00104# => romdata <= X"86A00003";
when 16#00105# => romdata <= X"84600002";
when 16#00106# => romdata <= X"C43FBFC8";
when 16#00107# => romdata <= X"C207BFF4";
when 16#00108# => romdata <= X"83286003";
when 16#00109# => romdata <= X"82078001";
when 16#0010A# => romdata <= X"C4187FC0";
when 16#0010B# => romdata <= X"84100003";
when 16#0010C# => romdata <= X"031FFFFF";
when 16#0010D# => romdata <= X"821063FF";
when 16#0010E# => romdata <= X"84088001";
when 16#0010F# => romdata <= X"C207A04C";
when 16#00110# => romdata <= X"C4204000";
when 16#00111# => romdata <= X"C207BFF4";
when 16#00112# => romdata <= X"82086001";
when 16#00113# => romdata <= X"84100001";
when 16#00114# => romdata <= X"C207A04C";
when 16#00115# => romdata <= X"8408A0FF";
when 16#00116# => romdata <= X"8528A01F";
when 16#00117# => romdata <= X"C8004000";
when 16#00118# => romdata <= X"071FFFFF";
when 16#00119# => romdata <= X"8610E3FF";
when 16#0011A# => romdata <= X"86090003";
when 16#0011B# => romdata <= X"8410C002";
when 16#0011C# => romdata <= X"C4204000";
when 16#0011D# => romdata <= X"81E80000";
when 16#0011E# => romdata <= X"81C3E008";
when 16#0011F# => romdata <= X"01000000";
when 16#00120# => romdata <= X"9DE3BF60";
when 16#00121# => romdata <= X"F027A044";
when 16#00122# => romdata <= X"F227A048";
when 16#00123# => romdata <= X"F427A04C";
when 16#00124# => romdata <= X"C207A044";
when 16#00125# => romdata <= X"C2004000";
when 16#00126# => romdata <= X"B4102000";
when 16#00127# => romdata <= X"B6100001";
when 16#00128# => romdata <= X"B8102000";
when 16#00129# => romdata <= X"3B1FFFFF";
when 16#0012A# => romdata <= X"BA1763FF";
when 16#0012B# => romdata <= X"B80E801C";
when 16#0012C# => romdata <= X"BA0EC01D";
when 16#0012D# => romdata <= X"F83FBFE0";
when 16#0012E# => romdata <= X"F81FBFE0";
when 16#0012F# => romdata <= X"BAA0001D";
when 16#00130# => romdata <= X"B860001C";
when 16#00131# => romdata <= X"F83FBFE8";
when 16#00132# => romdata <= X"C207A048";
when 16#00133# => romdata <= X"C2004000";
when 16#00134# => romdata <= X"B4102000";
when 16#00135# => romdata <= X"B6100001";
when 16#00136# => romdata <= X"B8102000";
when 16#00137# => romdata <= X"3B1FFFFF";
when 16#00138# => romdata <= X"BA1763FF";
when 16#00139# => romdata <= X"B80E801C";
when 16#0013A# => romdata <= X"BA0EC01D";
when 16#0013B# => romdata <= X"F83FBFD0";
when 16#0013C# => romdata <= X"F81FBFD0";
when 16#0013D# => romdata <= X"BAA0001D";
when 16#0013E# => romdata <= X"B860001C";
when 16#0013F# => romdata <= X"F83FBFD8";
when 16#00140# => romdata <= X"C207A044";
when 16#00141# => romdata <= X"C2004000";
when 16#00142# => romdata <= X"8330601F";
when 16#00143# => romdata <= X"820860FF";
when 16#00144# => romdata <= X"83286003";
when 16#00145# => romdata <= X"82078001";
when 16#00146# => romdata <= X"F4187FE0";
when 16#00147# => romdata <= X"C207A048";
when 16#00148# => romdata <= X"C2004000";
when 16#00149# => romdata <= X"8330601F";
when 16#0014A# => romdata <= X"820860FF";
when 16#0014B# => romdata <= X"83286003";
when 16#0014C# => romdata <= X"82078001";
when 16#0014D# => romdata <= X"F8187FD0";
when 16#0014E# => romdata <= X"BAA6C01D";
when 16#0014F# => romdata <= X"B866801C";
when 16#00150# => romdata <= X"F83FBFF8";
when 16#00151# => romdata <= X"F81FBFF8";
when 16#00152# => romdata <= X"8737201F";
when 16#00153# => romdata <= X"84102000";
when 16#00154# => romdata <= X"C627BFF4";
when 16#00155# => romdata <= X"C41FBFF8";
when 16#00156# => romdata <= X"C43FBFC0";
when 16#00157# => romdata <= X"C41FBFF8";
when 16#00158# => romdata <= X"86A00003";
when 16#00159# => romdata <= X"84600002";
when 16#0015A# => romdata <= X"C43FBFC8";
when 16#0015B# => romdata <= X"C207BFF4";
when 16#0015C# => romdata <= X"83286003";
when 16#0015D# => romdata <= X"82078001";
when 16#0015E# => romdata <= X"C4187FC0";
when 16#0015F# => romdata <= X"84100003";
when 16#00160# => romdata <= X"031FFFFF";
when 16#00161# => romdata <= X"821063FF";
when 16#00162# => romdata <= X"84088001";
when 16#00163# => romdata <= X"C207A04C";
when 16#00164# => romdata <= X"C4204000";
when 16#00165# => romdata <= X"C207BFF4";
when 16#00166# => romdata <= X"82086001";
when 16#00167# => romdata <= X"84100001";
when 16#00168# => romdata <= X"C207A04C";
when 16#00169# => romdata <= X"8408A0FF";
when 16#0016A# => romdata <= X"8528A01F";
when 16#0016B# => romdata <= X"C8004000";
when 16#0016C# => romdata <= X"071FFFFF";
when 16#0016D# => romdata <= X"8610E3FF";
when 16#0016E# => romdata <= X"86090003";
when 16#0016F# => romdata <= X"8410C002";
when 16#00170# => romdata <= X"C4204000";
when 16#00171# => romdata <= X"81E80000";
when 16#00172# => romdata <= X"81C3E008";
when 16#00173# => romdata <= X"01000000";
when 16#00174# => romdata <= X"9DE3BF98";
when 16#00175# => romdata <= X"F027A044";
when 16#00176# => romdata <= X"F227A048";
when 16#00177# => romdata <= X"8207BFFC";
when 16#00178# => romdata <= X"D007A044";
when 16#00179# => romdata <= X"D207A048";
when 16#0017A# => romdata <= X"94100001";
when 16#0017B# => romdata <= X"7FFFFFA5";
when 16#0017C# => romdata <= X"01000000";
when 16#0017D# => romdata <= X"C207BFFC";
when 16#0017E# => romdata <= X"80A06000";
when 16#0017F# => romdata <= X"12800005";
when 16#00180# => romdata <= X"01000000";
when 16#00181# => romdata <= X"82102000";
when 16#00182# => romdata <= X"1080000C";
when 16#00183# => romdata <= X"01000000";
when 16#00184# => romdata <= X"C407BFFC";
when 16#00185# => romdata <= X"03200000";
when 16#00186# => romdata <= X"82088001";
when 16#00187# => romdata <= X"80A06000";
when 16#00188# => romdata <= X"02800005";
when 16#00189# => romdata <= X"01000000";
when 16#0018A# => romdata <= X"82103FFF";
when 16#0018B# => romdata <= X"10800003";
when 16#0018C# => romdata <= X"01000000";
when 16#0018D# => romdata <= X"82102001";
when 16#0018E# => romdata <= X"B0100001";
when 16#0018F# => romdata <= X"81E80000";
when 16#00190# => romdata <= X"81C3E008";
when 16#00191# => romdata <= X"01000000";
when 16#00192# => romdata <= X"9DE3BFA0";
when 16#00193# => romdata <= X"F027A044";
when 16#00194# => romdata <= X"F227A048";
when 16#00195# => romdata <= X"C207A044";
when 16#00196# => romdata <= X"C4004000";
when 16#00197# => romdata <= X"C207A048";
when 16#00198# => romdata <= X"C4204000";
when 16#00199# => romdata <= X"C207A048";
when 16#0019A# => romdata <= X"C6004000";
when 16#0019B# => romdata <= X"051FFFFF";
when 16#0019C# => romdata <= X"8410A3FF";
when 16#0019D# => romdata <= X"8408C002";
when 16#0019E# => romdata <= X"C4204000";
when 16#0019F# => romdata <= X"81E80000";
when 16#001A0# => romdata <= X"81C3E008";
when 16#001A1# => romdata <= X"01000000";
when 16#001A2# => romdata <= X"9DE3BF98";
when 16#001A3# => romdata <= X"F027A044";
when 16#001A4# => romdata <= X"F227A048";
when 16#001A5# => romdata <= X"8207BFFC";
when 16#001A6# => romdata <= X"D007A044";
when 16#001A7# => romdata <= X"D207A048";
when 16#001A8# => romdata <= X"94100001";
when 16#001A9# => romdata <= X"7FFFFF77";
when 16#001AA# => romdata <= X"01000000";
when 16#001AB# => romdata <= X"C407BFFC";
when 16#001AC# => romdata <= X"03200000";
when 16#001AD# => romdata <= X"82088001";
when 16#001AE# => romdata <= X"82186000";
when 16#001AF# => romdata <= X"80A00001";
when 16#001B0# => romdata <= X"82603FFF";
when 16#001B1# => romdata <= X"820860FF";
when 16#001B2# => romdata <= X"B0100001";
when 16#001B3# => romdata <= X"81E80000";
when 16#001B4# => romdata <= X"81C3E008";
when 16#001B5# => romdata <= X"01000000";
when 16#001B6# => romdata <= X"9DE3BF98";
when 16#001B7# => romdata <= X"F027A044";
when 16#001B8# => romdata <= X"F227A048";
when 16#001B9# => romdata <= X"8207BFFC";
when 16#001BA# => romdata <= X"D007A048";
when 16#001BB# => romdata <= X"D207A044";
when 16#001BC# => romdata <= X"94100001";
when 16#001BD# => romdata <= X"7FFFFF63";
when 16#001BE# => romdata <= X"01000000";
when 16#001BF# => romdata <= X"C407BFFC";
when 16#001C0# => romdata <= X"03200000";
when 16#001C1# => romdata <= X"82088001";
when 16#001C2# => romdata <= X"82186000";
when 16#001C3# => romdata <= X"80A00001";
when 16#001C4# => romdata <= X"82603FFF";
when 16#001C5# => romdata <= X"820860FF";
when 16#001C6# => romdata <= X"B0100001";
when 16#001C7# => romdata <= X"81E80000";
when 16#001C8# => romdata <= X"81C3E008";
when 16#001C9# => romdata <= X"01000000";
when 16#001CA# => romdata <= X"9DE3BF98";
when 16#001CB# => romdata <= X"F027A044";
when 16#001CC# => romdata <= X"F227A048";
when 16#001CD# => romdata <= X"F427A04C";
when 16#001CE# => romdata <= X"C207A04C";
when 16#001CF# => romdata <= X"C407A044";
when 16#001D0# => romdata <= X"C400A034";
when 16#001D1# => romdata <= X"C4204000";
when 16#001D2# => romdata <= X"C027BFFC";
when 16#001D3# => romdata <= X"1080001A";
when 16#001D4# => romdata <= X"01000000";
when 16#001D5# => romdata <= X"C207BFFC";
when 16#001D6# => romdata <= X"83286002";
when 16#001D7# => romdata <= X"C407A044";
when 16#001D8# => romdata <= X"86008001";
when 16#001D9# => romdata <= X"C207BFFC";
when 16#001DA# => romdata <= X"83286002";
when 16#001DB# => romdata <= X"C407A048";
when 16#001DC# => romdata <= X"82008001";
when 16#001DD# => romdata <= X"C4004000";
when 16#001DE# => romdata <= X"8207BFF8";
when 16#001DF# => romdata <= X"90100003";
when 16#001E0# => romdata <= X"92100002";
when 16#001E1# => romdata <= X"94100001";
when 16#001E2# => romdata <= X"7FFFFEB2";
when 16#001E3# => romdata <= X"01000000";
when 16#001E4# => romdata <= X"8207BFF8";
when 16#001E5# => romdata <= X"D007A04C";
when 16#001E6# => romdata <= X"92100001";
when 16#001E7# => romdata <= X"D407A04C";
when 16#001E8# => romdata <= X"7FFFFEE4";
when 16#001E9# => romdata <= X"01000000";
when 16#001EA# => romdata <= X"C207BFFC";
when 16#001EB# => romdata <= X"82006001";
when 16#001EC# => romdata <= X"C227BFFC";
when 16#001ED# => romdata <= X"C207BFFC";
when 16#001EE# => romdata <= X"80A0600C";
when 16#001EF# => romdata <= X"04BFFFE6";
when 16#001F0# => romdata <= X"01000000";
when 16#001F1# => romdata <= X"81E80000";
when 16#001F2# => romdata <= X"81C3E008";
when 16#001F3# => romdata <= X"01000000";
when 16#001F4# => romdata <= X"9DE3BF68";
when 16#001F5# => romdata <= X"F027A044";
when 16#001F6# => romdata <= X"F227A048";
when 16#001F7# => romdata <= X"F427A04C";
when 16#001F8# => romdata <= X"F627A050";
when 16#001F9# => romdata <= X"C027BFFC";
when 16#001FA# => romdata <= X"1080000D";
when 16#001FB# => romdata <= X"01000000";
when 16#001FC# => romdata <= X"0310000B";
when 16#001FD# => romdata <= X"841062B8";
when 16#001FE# => romdata <= X"C207BFFC";
when 16#001FF# => romdata <= X"83286002";
when 16#00200# => romdata <= X"0710000A";
when 16#00201# => romdata <= X"8610E3A0";
when 16#00202# => romdata <= X"C600C000";
when 16#00203# => romdata <= X"C6208001";
when 16#00204# => romdata <= X"C207BFFC";
when 16#00205# => romdata <= X"82006001";
when 16#00206# => romdata <= X"C227BFFC";
when 16#00207# => romdata <= X"C207BFFC";
when 16#00208# => romdata <= X"80A06007";
when 16#00209# => romdata <= X"04BFFFF3";
when 16#0020A# => romdata <= X"01000000";
when 16#0020B# => romdata <= X"C027BFFC";
when 16#0020C# => romdata <= X"1080000F";
when 16#0020D# => romdata <= X"01000000";
when 16#0020E# => romdata <= X"C207BFFC";
when 16#0020F# => romdata <= X"82006008";
when 16#00210# => romdata <= X"C407BFFC";
when 16#00211# => romdata <= X"8528A002";
when 16#00212# => romdata <= X"C607A044";
when 16#00213# => romdata <= X"8600C002";
when 16#00214# => romdata <= X"05100009";
when 16#00215# => romdata <= X"8410A00C";
when 16#00216# => romdata <= X"83286002";
when 16#00217# => romdata <= X"C6208001";
when 16#00218# => romdata <= X"C207BFFC";
when 16#00219# => romdata <= X"82006001";
when 16#0021A# => romdata <= X"C227BFFC";
when 16#0021B# => romdata <= X"C207BFFC";
when 16#0021C# => romdata <= X"80A06002";
when 16#0021D# => romdata <= X"04BFFFF1";
when 16#0021E# => romdata <= X"01000000";
when 16#0021F# => romdata <= X"03100009";
when 16#00220# => romdata <= X"8210600C";
when 16#00221# => romdata <= X"C407A04C";
when 16#00222# => romdata <= X"C420602C";
when 16#00223# => romdata <= X"03100009";
when 16#00224# => romdata <= X"8210600C";
when 16#00225# => romdata <= X"C407A048";
when 16#00226# => romdata <= X"C4206030";
when 16#00227# => romdata <= X"C027BFFC";
when 16#00228# => romdata <= X"10800074";
when 16#00229# => romdata <= X"01000000";
when 16#0022A# => romdata <= X"C027BFF8";
when 16#0022B# => romdata <= X"1080000E";
when 16#0022C# => romdata <= X"01000000";
when 16#0022D# => romdata <= X"C207BFF8";
when 16#0022E# => romdata <= X"83286002";
when 16#0022F# => romdata <= X"82078001";
when 16#00230# => romdata <= X"0510000B";
when 16#00231# => romdata <= X"8610A2B8";
when 16#00232# => romdata <= X"C407BFF8";
when 16#00233# => romdata <= X"8528A002";
when 16#00234# => romdata <= X"C400C002";
when 16#00235# => romdata <= X"C4207FD8";
when 16#00236# => romdata <= X"C207BFF8";
when 16#00237# => romdata <= X"82006001";
when 16#00238# => romdata <= X"C227BFF8";
when 16#00239# => romdata <= X"C207BFF8";
when 16#0023A# => romdata <= X"80A06007";
when 16#0023B# => romdata <= X"04BFFFF2";
when 16#0023C# => romdata <= X"01000000";
when 16#0023D# => romdata <= X"C027BFF8";
when 16#0023E# => romdata <= X"1080001F";
when 16#0023F# => romdata <= X"01000000";
when 16#00240# => romdata <= X"C207BFF8";
when 16#00241# => romdata <= X"83286003";
when 16#00242# => romdata <= X"85286003";
when 16#00243# => romdata <= X"84208001";
when 16#00244# => romdata <= X"03100009";
when 16#00245# => romdata <= X"82106040";
when 16#00246# => romdata <= X"84008001";
when 16#00247# => romdata <= X"8207BFD4";
when 16#00248# => romdata <= X"90100002";
when 16#00249# => romdata <= X"05100009";
when 16#0024A# => romdata <= X"9210A00C";
when 16#0024B# => romdata <= X"94100001";
when 16#0024C# => romdata <= X"7FFFFF7E";
when 16#0024D# => romdata <= X"01000000";
when 16#0024E# => romdata <= X"C407BFD4";
when 16#0024F# => romdata <= X"03200000";
when 16#00250# => romdata <= X"82088001";
when 16#00251# => romdata <= X"80A06000";
when 16#00252# => romdata <= X"12800008";
when 16#00253# => romdata <= X"01000000";
when 16#00254# => romdata <= X"0310000B";
when 16#00255# => romdata <= X"841062B8";
when 16#00256# => romdata <= X"C207BFF8";
when 16#00257# => romdata <= X"83286002";
when 16#00258# => romdata <= X"C607BFD4";
when 16#00259# => romdata <= X"C6208001";
when 16#0025A# => romdata <= X"C207BFF8";
when 16#0025B# => romdata <= X"82006001";
when 16#0025C# => romdata <= X"C227BFF8";
when 16#0025D# => romdata <= X"C207BFF8";
when 16#0025E# => romdata <= X"80A06007";
when 16#0025F# => romdata <= X"04BFFFE1";
when 16#00260# => romdata <= X"01000000";
when 16#00261# => romdata <= X"0310000A";
when 16#00262# => romdata <= X"821063A0";
when 16#00263# => romdata <= X"C2004000";
when 16#00264# => romdata <= X"C227BFD0";
when 16#00265# => romdata <= X"C027BFC8";
when 16#00266# => romdata <= X"82102015";
when 16#00267# => romdata <= X"C237BFCA";
when 16#00268# => romdata <= X"C027BFF8";
when 16#00269# => romdata <= X"10800021";
when 16#0026A# => romdata <= X"01000000";
when 16#0026B# => romdata <= X"C207BFF8";
when 16#0026C# => romdata <= X"85286002";
when 16#0026D# => romdata <= X"0310000B";
when 16#0026E# => romdata <= X"821062B8";
when 16#0026F# => romdata <= X"86008001";
when 16#00270# => romdata <= X"C207BFF8";
when 16#00271# => romdata <= X"83286002";
when 16#00272# => romdata <= X"8407BFD8";
when 16#00273# => romdata <= X"84008001";
when 16#00274# => romdata <= X"8207BFCC";
when 16#00275# => romdata <= X"90100003";
when 16#00276# => romdata <= X"92100002";
when 16#00277# => romdata <= X"94100001";
when 16#00278# => romdata <= X"7FFFFEA8";
when 16#00279# => romdata <= X"01000000";
when 16#0027A# => romdata <= X"C407BFCC";
when 16#0027B# => romdata <= X"031FFFFF";
when 16#0027C# => romdata <= X"821063FF";
when 16#0027D# => romdata <= X"82088001";
when 16#0027E# => romdata <= X"C227BFCC";
when 16#0027F# => romdata <= X"8607BFD0";
when 16#00280# => romdata <= X"8407BFCC";
when 16#00281# => romdata <= X"8207BFD0";
when 16#00282# => romdata <= X"90100003";
when 16#00283# => romdata <= X"92100002";
when 16#00284# => romdata <= X"94100001";
when 16#00285# => romdata <= X"7FFFFE47";
when 16#00286# => romdata <= X"01000000";
when 16#00287# => romdata <= X"C207BFF8";
when 16#00288# => romdata <= X"82006001";
when 16#00289# => romdata <= X"C227BFF8";
when 16#0028A# => romdata <= X"C207BFF8";
when 16#0028B# => romdata <= X"80A06007";
when 16#0028C# => romdata <= X"04BFFFDF";
when 16#0028D# => romdata <= X"01000000";
when 16#0028E# => romdata <= X"8407BFD0";
when 16#0028F# => romdata <= X"8207BFC8";
when 16#00290# => romdata <= X"90100002";
when 16#00291# => romdata <= X"92100001";
when 16#00292# => romdata <= X"7FFFFF24";
when 16#00293# => romdata <= X"01000000";
when 16#00294# => romdata <= X"82100008";
when 16#00295# => romdata <= X"820860FF";
when 16#00296# => romdata <= X"80A06000";
when 16#00297# => romdata <= X"1280000B";
when 16#00298# => romdata <= X"01000000";
when 16#00299# => romdata <= X"C207BFFC";
when 16#0029A# => romdata <= X"82006001";
when 16#0029B# => romdata <= X"C227BFFC";
when 16#0029C# => romdata <= X"C207BFFC";
when 16#0029D# => romdata <= X"80A06018";
when 16#0029E# => romdata <= X"04BFFF8C";
when 16#0029F# => romdata <= X"01000000";
when 16#002A0# => romdata <= X"10800003";
when 16#002A1# => romdata <= X"01000000";
when 16#002A2# => romdata <= X"01000000";
when 16#002A3# => romdata <= X"03100009";
when 16#002A4# => romdata <= X"90106200";
when 16#002A5# => romdata <= X"03100009";
when 16#002A6# => romdata <= X"9210600C";
when 16#002A7# => romdata <= X"D407A050";
when 16#002A8# => romdata <= X"7FFFFF22";
when 16#002A9# => romdata <= X"01000000";
when 16#002AA# => romdata <= X"C027BFFC";
when 16#002AB# => romdata <= X"C207BFFC";
when 16#002AC# => romdata <= X"82006001";
when 16#002AD# => romdata <= X"C227BFFC";
when 16#002AE# => romdata <= X"C207BFFC";
when 16#002AF# => romdata <= X"82006001";
when 16#002B0# => romdata <= X"C227BFFC";
when 16#002B1# => romdata <= X"C207BFFC";
when 16#002B2# => romdata <= X"82006001";
when 16#002B3# => romdata <= X"C227BFFC";
when 16#002B4# => romdata <= X"C207BFFC";
when 16#002B5# => romdata <= X"82006001";
when 16#002B6# => romdata <= X"C227BFFC";
when 16#002B7# => romdata <= X"C207BFFC";
when 16#002B8# => romdata <= X"82006001";
when 16#002B9# => romdata <= X"C227BFFC";
when 16#002BA# => romdata <= X"C207BFFC";
when 16#002BB# => romdata <= X"82006001";
when 16#002BC# => romdata <= X"C227BFFC";
when 16#002BD# => romdata <= X"C207BFFC";
when 16#002BE# => romdata <= X"82006001";
when 16#002BF# => romdata <= X"C227BFFC";
when 16#002C0# => romdata <= X"C207BFFC";
when 16#002C1# => romdata <= X"82006001";
when 16#002C2# => romdata <= X"C227BFFC";
when 16#002C3# => romdata <= X"81E80000";
when 16#002C4# => romdata <= X"81C3E008";
when 16#002C5# => romdata <= X"01000000";
when 16#002C6# => romdata <= X"9DE3BFA0";
when 16#002C7# => romdata <= X"82100018";
when 16#002C8# => romdata <= X"C237A044";
when 16#002C9# => romdata <= X"03100009";
when 16#002CA# => romdata <= X"82106238";
when 16#002CB# => romdata <= X"C417A044";
when 16#002CC# => romdata <= X"C4304000";
when 16#002CD# => romdata <= X"81E80000";
when 16#002CE# => romdata <= X"81C3E008";
when 16#002CF# => romdata <= X"01000000";
when 16#002D0# => romdata <= X"9DE3BF98";
when 16#002D1# => romdata <= X"03100009";
when 16#002D2# => romdata <= X"82106238";
when 16#002D3# => romdata <= X"C2104000";
when 16#002D4# => romdata <= X"83286010";
when 16#002D5# => romdata <= X"83306010";
when 16#002D6# => romdata <= X"83306002";
when 16#002D7# => romdata <= X"84100001";
when 16#002D8# => romdata <= X"03100009";
when 16#002D9# => romdata <= X"82106238";
when 16#002DA# => romdata <= X"C2104000";
when 16#002DB# => romdata <= X"82188001";
when 16#002DC# => romdata <= X"84100001";
when 16#002DD# => romdata <= X"03100009";
when 16#002DE# => romdata <= X"82106238";
when 16#002DF# => romdata <= X"C2104000";
when 16#002E0# => romdata <= X"83286010";
when 16#002E1# => romdata <= X"83306010";
when 16#002E2# => romdata <= X"83306003";
when 16#002E3# => romdata <= X"82188001";
when 16#002E4# => romdata <= X"84100001";
when 16#002E5# => romdata <= X"03100009";
when 16#002E6# => romdata <= X"82106238";
when 16#002E7# => romdata <= X"C2104000";
when 16#002E8# => romdata <= X"83286010";
when 16#002E9# => romdata <= X"83306010";
when 16#002EA# => romdata <= X"83306005";
when 16#002EB# => romdata <= X"82188001";
when 16#002EC# => romdata <= X"82086001";
when 16#002ED# => romdata <= X"C237BFFE";
when 16#002EE# => romdata <= X"03100009";
when 16#002EF# => romdata <= X"82106238";
when 16#002F0# => romdata <= X"C2104000";
when 16#002F1# => romdata <= X"83286010";
when 16#002F2# => romdata <= X"83306010";
when 16#002F3# => romdata <= X"83306001";
when 16#002F4# => romdata <= X"84100001";
when 16#002F5# => romdata <= X"C217BFFE";
when 16#002F6# => romdata <= X"83286010";
when 16#002F7# => romdata <= X"83306010";
when 16#002F8# => romdata <= X"8328600F";
when 16#002F9# => romdata <= X"82108001";
when 16#002FA# => romdata <= X"84100001";
when 16#002FB# => romdata <= X"03100009";
when 16#002FC# => romdata <= X"82106238";
when 16#002FD# => romdata <= X"C4304000";
when 16#002FE# => romdata <= X"03100009";
when 16#002FF# => romdata <= X"82106238";
when 16#00300# => romdata <= X"C2104000";
when 16#00301# => romdata <= X"83286010";
when 16#00302# => romdata <= X"83306010";
when 16#00303# => romdata <= X"B0100001";
when 16#00304# => romdata <= X"81E80000";
when 16#00305# => romdata <= X"81C3E008";
when 16#00306# => romdata <= X"01000000";
when 16#00307# => romdata <= X"9DE3BF88";
when 16#00308# => romdata <= X"F027A044";
when 16#00309# => romdata <= X"82102001";
when 16#0030A# => romdata <= X"C227BFFC";
when 16#0030B# => romdata <= X"C027BFF8";
when 16#0030C# => romdata <= X"10800038";
when 16#0030D# => romdata <= X"01000000";
when 16#0030E# => romdata <= X"C027BFFC";
when 16#0030F# => romdata <= X"C027BFF4";
when 16#00310# => romdata <= X"1080002A";
when 16#00311# => romdata <= X"01000000";
when 16#00312# => romdata <= X"C207BFF4";
when 16#00313# => romdata <= X"82006001";
when 16#00314# => romdata <= X"C227BFF0";
when 16#00315# => romdata <= X"C207BFF4";
when 16#00316# => romdata <= X"C407A044";
when 16#00317# => romdata <= X"82008001";
when 16#00318# => romdata <= X"C4084000";
when 16#00319# => romdata <= X"C207BFF0";
when 16#0031A# => romdata <= X"C607A044";
when 16#0031B# => romdata <= X"8200C001";
when 16#0031C# => romdata <= X"C2084000";
when 16#0031D# => romdata <= X"8408A0FF";
when 16#0031E# => romdata <= X"820860FF";
when 16#0031F# => romdata <= X"80A08001";
when 16#00320# => romdata <= X"08800017";
when 16#00321# => romdata <= X"01000000";
when 16#00322# => romdata <= X"C207BFF4";
when 16#00323# => romdata <= X"C407A044";
when 16#00324# => romdata <= X"82008001";
when 16#00325# => romdata <= X"C2084000";
when 16#00326# => romdata <= X"820860FF";
when 16#00327# => romdata <= X"C227BFEC";
when 16#00328# => romdata <= X"C207BFF4";
when 16#00329# => romdata <= X"C407A044";
when 16#0032A# => romdata <= X"82008001";
when 16#0032B# => romdata <= X"C407BFF0";
when 16#0032C# => romdata <= X"C607A044";
when 16#0032D# => romdata <= X"8400C002";
when 16#0032E# => romdata <= X"C4088000";
when 16#0032F# => romdata <= X"C4284000";
when 16#00330# => romdata <= X"C207BFF0";
when 16#00331# => romdata <= X"C407A044";
when 16#00332# => romdata <= X"82008001";
when 16#00333# => romdata <= X"C407BFEC";
when 16#00334# => romdata <= X"C4284000";
when 16#00335# => romdata <= X"82102001";
when 16#00336# => romdata <= X"C227BFFC";
when 16#00337# => romdata <= X"C207BFF4";
when 16#00338# => romdata <= X"82006001";
when 16#00339# => romdata <= X"C227BFF4";
when 16#0033A# => romdata <= X"84102013";
when 16#0033B# => romdata <= X"C207BFF8";
when 16#0033C# => romdata <= X"84208001";
when 16#0033D# => romdata <= X"C207BFF4";
when 16#0033E# => romdata <= X"80A08001";
when 16#0033F# => romdata <= X"14BFFFD3";
when 16#00340# => romdata <= X"01000000";
when 16#00341# => romdata <= X"C207BFF8";
when 16#00342# => romdata <= X"82006001";
when 16#00343# => romdata <= X"C227BFF8";
when 16#00344# => romdata <= X"C207BFF8";
when 16#00345# => romdata <= X"80A06013";
when 16#00346# => romdata <= X"14800006";
when 16#00347# => romdata <= X"01000000";
when 16#00348# => romdata <= X"C207BFFC";
when 16#00349# => romdata <= X"80A06000";
when 16#0034A# => romdata <= X"12BFFFC4";
when 16#0034B# => romdata <= X"01000000";
when 16#0034C# => romdata <= X"81E80000";
when 16#0034D# => romdata <= X"81C3E008";
when 16#0034E# => romdata <= X"01000000";
when 16#0034F# => romdata <= X"9DE3BF98";
when 16#00350# => romdata <= X"BB444000";
when 16#00351# => romdata <= X"FA27BFFC";
when 16#00352# => romdata <= X"C207BFFC";
when 16#00353# => romdata <= X"B0100001";
when 16#00354# => romdata <= X"81E80000";
when 16#00355# => romdata <= X"81C3E008";
when 16#00356# => romdata <= X"01000000";
when 16#00357# => romdata <= X"9DE3BFA0";
when 16#00358# => romdata <= X"7FFFFFF7";
when 16#00359# => romdata <= X"01000000";
when 16#0035A# => romdata <= X"82100008";
when 16#0035B# => romdata <= X"8330601C";
when 16#0035C# => romdata <= X"B0100001";
when 16#0035D# => romdata <= X"81E80000";
when 16#0035E# => romdata <= X"81C3E008";
when 16#0035F# => romdata <= X"01000000";
when 16#00360# => romdata <= X"9DE3BFA0";
when 16#00361# => romdata <= X"F027A044";
when 16#00362# => romdata <= X"C207A044";
when 16#00363# => romdata <= X"8208600F";
when 16#00364# => romdata <= X"C227A044";
when 16#00365# => romdata <= X"03200000";
when 16#00366# => romdata <= X"82106210";
when 16#00367# => romdata <= X"05200000";
when 16#00368# => romdata <= X"8410A210";
when 16#00369# => romdata <= X"C6008000";
when 16#0036A# => romdata <= X"88102001";
when 16#0036B# => romdata <= X"C407A044";
when 16#0036C# => romdata <= X"85290002";
when 16#0036D# => romdata <= X"8410C002";
when 16#0036E# => romdata <= X"C4204000";
when 16#0036F# => romdata <= X"81E80000";
when 16#00370# => romdata <= X"81C3E008";
when 16#00371# => romdata <= X"01000000";
when 16#00372# => romdata <= X"9DE3BFA0";
when 16#00373# => romdata <= X"F027A044";
when 16#00374# => romdata <= X"C207A044";
when 16#00375# => romdata <= X"8208600F";
when 16#00376# => romdata <= X"C227A044";
when 16#00377# => romdata <= X"03200000";
when 16#00378# => romdata <= X"82106210";
when 16#00379# => romdata <= X"05200000";
when 16#0037A# => romdata <= X"8410A210";
when 16#0037B# => romdata <= X"C6008000";
when 16#0037C# => romdata <= X"88102001";
when 16#0037D# => romdata <= X"C407A044";
when 16#0037E# => romdata <= X"85290002";
when 16#0037F# => romdata <= X"84380002";
when 16#00380# => romdata <= X"8408C002";
when 16#00381# => romdata <= X"C4204000";
when 16#00382# => romdata <= X"81E80000";
when 16#00383# => romdata <= X"81C3E008";
when 16#00384# => romdata <= X"01000000";
when 16#00385# => romdata <= X"9DE3BF98";
when 16#00386# => romdata <= X"F027A044";
when 16#00387# => romdata <= X"7FFFFF49";
when 16#00388# => romdata <= X"01000000";
when 16#00389# => romdata <= X"82100008";
when 16#0038A# => romdata <= X"83286010";
when 16#0038B# => romdata <= X"83306010";
when 16#0038C# => romdata <= X"C227BFFC";
when 16#0038D# => romdata <= X"C207BFFC";
when 16#0038E# => romdata <= X"82086001";
when 16#0038F# => romdata <= X"C227BFF8";
when 16#00390# => romdata <= X"C207BFFC";
when 16#00391# => romdata <= X"83286003";
when 16#00392# => romdata <= X"C227BFFC";
when 16#00393# => romdata <= X"C207A044";
when 16#00394# => romdata <= X"C407BFFC";
when 16#00395# => romdata <= X"C4204000";
when 16#00396# => romdata <= X"C207BFF8";
when 16#00397# => romdata <= X"82086001";
when 16#00398# => romdata <= X"84100001";
when 16#00399# => romdata <= X"C207A044";
when 16#0039A# => romdata <= X"8408A0FF";
when 16#0039B# => romdata <= X"8528A01F";
when 16#0039C# => romdata <= X"C8004000";
when 16#0039D# => romdata <= X"071FFFFF";
when 16#0039E# => romdata <= X"8610E3FF";
when 16#0039F# => romdata <= X"86090003";
when 16#003A0# => romdata <= X"8410C002";
when 16#003A1# => romdata <= X"C4204000";
when 16#003A2# => romdata <= X"81E80000";
when 16#003A3# => romdata <= X"81C3E008";
when 16#003A4# => romdata <= X"01000000";
when 16#003A5# => romdata <= X"9DE3BF98";
when 16#003A6# => romdata <= X"F027A044";
when 16#003A7# => romdata <= X"7FFFFF29";
when 16#003A8# => romdata <= X"01000000";
when 16#003A9# => romdata <= X"82100008";
when 16#003AA# => romdata <= X"83286010";
when 16#003AB# => romdata <= X"83306010";
when 16#003AC# => romdata <= X"C227BFFC";
when 16#003AD# => romdata <= X"C207BFFC";
when 16#003AE# => romdata <= X"82086001";
when 16#003AF# => romdata <= X"C227BFF8";
when 16#003B0# => romdata <= X"C207BFFC";
when 16#003B1# => romdata <= X"83286001";
when 16#003B2# => romdata <= X"C227BFFC";
when 16#003B3# => romdata <= X"C207A044";
when 16#003B4# => romdata <= X"C407BFFC";
when 16#003B5# => romdata <= X"C4204000";
when 16#003B6# => romdata <= X"C207BFF8";
when 16#003B7# => romdata <= X"82086001";
when 16#003B8# => romdata <= X"84100001";
when 16#003B9# => romdata <= X"C207A044";
when 16#003BA# => romdata <= X"8408A0FF";
when 16#003BB# => romdata <= X"8528A01F";
when 16#003BC# => romdata <= X"C8004000";
when 16#003BD# => romdata <= X"071FFFFF";
when 16#003BE# => romdata <= X"8610E3FF";
when 16#003BF# => romdata <= X"86090003";
when 16#003C0# => romdata <= X"8410C002";
when 16#003C1# => romdata <= X"C4204000";
when 16#003C2# => romdata <= X"81E80000";
when 16#003C3# => romdata <= X"81C3E008";
when 16#003C4# => romdata <= X"01000000";
when 16#003C5# => romdata <= X"9DE3BF70";
when 16#003C6# => romdata <= X"7FFFFF91";
when 16#003C7# => romdata <= X"01000000";
when 16#003C8# => romdata <= X"82100008";
when 16#003C9# => romdata <= X"80A06000";
when 16#003CA# => romdata <= X"1280007D";
when 16#003CB# => romdata <= X"01000000";
when 16#003CC# => romdata <= X"03100009";
when 16#003CD# => romdata <= X"82106240";
when 16#003CE# => romdata <= X"84102001";
when 16#003CF# => romdata <= X"C4284000";
when 16#003D0# => romdata <= X"03100009";
when 16#003D1# => romdata <= X"82106240";
when 16#003D2# => romdata <= X"84102001";
when 16#003D3# => romdata <= X"C4284000";
when 16#003D4# => romdata <= X"C027BFE0";
when 16#003D5# => romdata <= X"C027BFE4";
when 16#003D6# => romdata <= X"C027BFE8";
when 16#003D7# => romdata <= X"0310000A";
when 16#003D8# => romdata <= X"821063A0";
when 16#003D9# => romdata <= X"C2004000";
when 16#003DA# => romdata <= X"C227BFE0";
when 16#003DB# => romdata <= X"0310000A";
when 16#003DC# => romdata <= X"821063A0";
when 16#003DD# => romdata <= X"C2004000";
when 16#003DE# => romdata <= X"C227BFE4";
when 16#003DF# => romdata <= X"0310000A";
when 16#003E0# => romdata <= X"821063A0";
when 16#003E1# => romdata <= X"C2004000";
when 16#003E2# => romdata <= X"C227BFE8";
when 16#003E3# => romdata <= X"0310000A";
when 16#003E4# => romdata <= X"821063A0";
when 16#003E5# => romdata <= X"C2004000";
when 16#003E6# => romdata <= X"C227BFD8";
when 16#003E7# => romdata <= X"01000000";
when 16#003E8# => romdata <= X"03100009";
when 16#003E9# => romdata <= X"8210623C";
when 16#003EA# => romdata <= X"C2004000";
when 16#003EB# => romdata <= X"C4004000";
when 16#003EC# => romdata <= X"03200000";
when 16#003ED# => romdata <= X"80A08001";
when 16#003EE# => romdata <= X"12BFFFFA";
when 16#003EF# => romdata <= X"01000000";
when 16#003F0# => romdata <= X"03100009";
when 16#003F1# => romdata <= X"8210623C";
when 16#003F2# => romdata <= X"C2004000";
when 16#003F3# => romdata <= X"C2006004";
when 16#003F4# => romdata <= X"C227BFDC";
when 16#003F5# => romdata <= X"03100009";
when 16#003F6# => romdata <= X"8210623C";
when 16#003F7# => romdata <= X"C2004000";
when 16#003F8# => romdata <= X"82006008";
when 16#003F9# => romdata <= X"C2004000";
when 16#003FA# => romdata <= X"C227BFF0";
when 16#003FB# => romdata <= X"03100009";
when 16#003FC# => romdata <= X"8210623C";
when 16#003FD# => romdata <= X"C2004000";
when 16#003FE# => romdata <= X"8200600C";
when 16#003FF# => romdata <= X"C2004000";
when 16#00400# => romdata <= X"83286010";
when 16#00401# => romdata <= X"83306010";
when 16#00402# => romdata <= X"90100001";
when 16#00403# => romdata <= X"7FFFFEC3";
when 16#00404# => romdata <= X"01000000";
when 16#00405# => romdata <= X"7FFFFECB";
when 16#00406# => romdata <= X"01000000";
when 16#00407# => romdata <= X"03100009";
when 16#00408# => romdata <= X"8210623C";
when 16#00409# => romdata <= X"C2004000";
when 16#0040A# => romdata <= X"82006010";
when 16#0040B# => romdata <= X"C2004000";
when 16#0040C# => romdata <= X"80A06000";
when 16#0040D# => romdata <= X"02800005";
when 16#0040E# => romdata <= X"01000000";
when 16#0040F# => romdata <= X"90102001";
when 16#00410# => romdata <= X"7FFFFF50";
when 16#00411# => romdata <= X"01000000";
when 16#00412# => romdata <= X"01000000";
when 16#00413# => romdata <= X"01000000";
when 16#00414# => romdata <= X"C027BFFC";
when 16#00415# => romdata <= X"10800025";
when 16#00416# => romdata <= X"01000000";
when 16#00417# => romdata <= X"8807BFE0";
when 16#00418# => romdata <= X"8607BFD8";
when 16#00419# => romdata <= X"8407BFDC";
when 16#0041A# => romdata <= X"8207BFD4";
when 16#0041B# => romdata <= X"90100004";
when 16#0041C# => romdata <= X"92100003";
when 16#0041D# => romdata <= X"94100002";
when 16#0041E# => romdata <= X"96100001";
when 16#0041F# => romdata <= X"7FFFFDD5";
when 16#00420# => romdata <= X"01000000";
when 16#00421# => romdata <= X"8207BFDC";
when 16#00422# => romdata <= X"90100001";
when 16#00423# => romdata <= X"7FFFFF62";
when 16#00424# => romdata <= X"01000000";
when 16#00425# => romdata <= X"8207BFD8";
when 16#00426# => romdata <= X"90100001";
when 16#00427# => romdata <= X"7FFFFF7E";
when 16#00428# => romdata <= X"01000000";
when 16#00429# => romdata <= X"8207BFE0";
when 16#0042A# => romdata <= X"90100001";
when 16#0042B# => romdata <= X"7FFFFF5A";
when 16#0042C# => romdata <= X"01000000";
when 16#0042D# => romdata <= X"8207BFE0";
when 16#0042E# => romdata <= X"82006004";
when 16#0042F# => romdata <= X"90100001";
when 16#00430# => romdata <= X"7FFFFF55";
when 16#00431# => romdata <= X"01000000";
when 16#00432# => romdata <= X"8207BFE0";
when 16#00433# => romdata <= X"82006008";
when 16#00434# => romdata <= X"90100001";
when 16#00435# => romdata <= X"7FFFFF50";
when 16#00436# => romdata <= X"01000000";
when 16#00437# => romdata <= X"C207BFFC";
when 16#00438# => romdata <= X"82006001";
when 16#00439# => romdata <= X"C227BFFC";
when 16#0043A# => romdata <= X"C407BFFC";
when 16#0043B# => romdata <= X"C207BFF0";
when 16#0043C# => romdata <= X"80A08001";
when 16#0043D# => romdata <= X"06BFFFDA";
when 16#0043E# => romdata <= X"01000000";
when 16#0043F# => romdata <= X"03100009";
when 16#00440# => romdata <= X"82106240";
when 16#00441# => romdata <= X"C0284000";
when 16#00442# => romdata <= X"03100009";
when 16#00443# => romdata <= X"82106240";
when 16#00444# => romdata <= X"C0284000";
when 16#00445# => romdata <= X"10800050";
when 16#00446# => romdata <= X"01000000";
when 16#00447# => romdata <= X"03100009";
when 16#00448# => romdata <= X"8210623C";
when 16#00449# => romdata <= X"C2004000";
when 16#0044A# => romdata <= X"8200600C";
when 16#0044B# => romdata <= X"C2004000";
when 16#0044C# => romdata <= X"C237BFF6";
when 16#0044D# => romdata <= X"0310000A";
when 16#0044E# => romdata <= X"821063A4";
when 16#0044F# => romdata <= X"C0204000";
when 16#00450# => romdata <= X"1080003E";
when 16#00451# => romdata <= X"01000000";
when 16#00452# => romdata <= X"C027BFF8";
when 16#00453# => romdata <= X"1080002C";
when 16#00454# => romdata <= X"01000000";
when 16#00455# => romdata <= X"C217BFF6";
when 16#00456# => romdata <= X"83286010";
when 16#00457# => romdata <= X"83306010";
when 16#00458# => romdata <= X"83306002";
when 16#00459# => romdata <= X"84100001";
when 16#0045A# => romdata <= X"C217BFF6";
when 16#0045B# => romdata <= X"82188001";
when 16#0045C# => romdata <= X"84100001";
when 16#0045D# => romdata <= X"C217BFF6";
when 16#0045E# => romdata <= X"83286010";
when 16#0045F# => romdata <= X"83306010";
when 16#00460# => romdata <= X"83306003";
when 16#00461# => romdata <= X"82188001";
when 16#00462# => romdata <= X"84100001";
when 16#00463# => romdata <= X"C217BFF6";
when 16#00464# => romdata <= X"83286010";
when 16#00465# => romdata <= X"83306010";
when 16#00466# => romdata <= X"83306005";
when 16#00467# => romdata <= X"82188001";
when 16#00468# => romdata <= X"82086001";
when 16#00469# => romdata <= X"C237BFEE";
when 16#0046A# => romdata <= X"C217BFF6";
when 16#0046B# => romdata <= X"83286010";
when 16#0046C# => romdata <= X"83306010";
when 16#0046D# => romdata <= X"83306001";
when 16#0046E# => romdata <= X"84100001";
when 16#0046F# => romdata <= X"C217BFEE";
when 16#00470# => romdata <= X"83286010";
when 16#00471# => romdata <= X"83306010";
when 16#00472# => romdata <= X"8328600F";
when 16#00473# => romdata <= X"82108001";
when 16#00474# => romdata <= X"C237BFF6";
when 16#00475# => romdata <= X"C217BFF6";
when 16#00476# => romdata <= X"84100001";
when 16#00477# => romdata <= X"0310000B";
when 16#00478# => romdata <= X"861062D8";
when 16#00479# => romdata <= X"C207BFF8";
when 16#0047A# => romdata <= X"8200C001";
when 16#0047B# => romdata <= X"C4284000";
when 16#0047C# => romdata <= X"C207BFF8";
when 16#0047D# => romdata <= X"82006001";
when 16#0047E# => romdata <= X"C227BFF8";
when 16#0047F# => romdata <= X"C207BFF8";
when 16#00480# => romdata <= X"80A06013";
when 16#00481# => romdata <= X"04BFFFD4";
when 16#00482# => romdata <= X"01000000";
when 16#00483# => romdata <= X"0310000B";
when 16#00484# => romdata <= X"901062D8";
when 16#00485# => romdata <= X"7FFFFE82";
when 16#00486# => romdata <= X"01000000";
when 16#00487# => romdata <= X"0310000A";
when 16#00488# => romdata <= X"821063A4";
when 16#00489# => romdata <= X"C2004000";
when 16#0048A# => romdata <= X"84006001";
when 16#0048B# => romdata <= X"0310000A";
when 16#0048C# => romdata <= X"821063A4";
when 16#0048D# => romdata <= X"C4204000";
when 16#0048E# => romdata <= X"03100009";
when 16#0048F# => romdata <= X"82106240";
when 16#00490# => romdata <= X"C2084000";
when 16#00491# => romdata <= X"820860FF";
when 16#00492# => romdata <= X"80A06001";
when 16#00493# => romdata <= X"02BFFFBF";
when 16#00494# => romdata <= X"01000000";
when 16#00495# => romdata <= X"B0100001";
when 16#00496# => romdata <= X"81E80000";
when 16#00497# => romdata <= X"81C3E008";
when 16#00498# => romdata <= X"01000000";
when 16#00499# => romdata <= X"92100008";
when 16#0049A# => romdata <= X"94102000";
when 16#0049B# => romdata <= X"90102000";
when 16#0049C# => romdata <= X"96102000";
when 16#0049D# => romdata <= X"8213C000";
when 16#0049E# => romdata <= X"40000002";
when 16#0049F# => romdata <= X"9E104000";
when 16#004A0# => romdata <= X"9DE3BFA0";
when 16#004A1# => romdata <= X"03100008";
when 16#004A2# => romdata <= X"FA006270";
when 16#004A3# => romdata <= X"D0076148";
when 16#004A4# => romdata <= X"80A22000";
when 16#004A5# => romdata <= X"02800034";
when 16#004A6# => romdata <= X"B8100018";
when 16#004A7# => romdata <= X"C2022004";
when 16#004A8# => romdata <= X"80A0601F";
when 16#004A9# => romdata <= X"04800015";
when 16#004AA# => romdata <= X"80A72000";
when 16#004AB# => romdata <= X"03000000";
when 16#004AC# => romdata <= X"82106000";
when 16#004AD# => romdata <= X"80A06000";
when 16#004AE# => romdata <= X"12800004";
when 16#004AF# => romdata <= X"B0103FFF";
when 16#004B0# => romdata <= X"81C7E008";
when 16#004B1# => romdata <= X"81E80000";
when 16#004B2# => romdata <= X"6FFFFB4E";
when 16#004B3# => romdata <= X"90102190";
when 16#004B4# => romdata <= X"80A22000";
when 16#004B5# => romdata <= X"02BFFFFB";
when 16#004B6# => romdata <= X"80A72000";
when 16#004B7# => romdata <= X"C2076148";
when 16#004B8# => romdata <= X"C2220000";
when 16#004B9# => romdata <= X"C0222004";
when 16#004BA# => romdata <= X"D0276148";
when 16#004BB# => romdata <= X"C0222188";
when 16#004BC# => romdata <= X"C022218C";
when 16#004BD# => romdata <= X"82102000";
when 16#004BE# => romdata <= X"02800011";
when 16#004BF# => romdata <= X"84006002";
when 16#004C0# => romdata <= X"C8022188";
when 16#004C1# => romdata <= X"BB286002";
when 16#004C2# => romdata <= X"84102001";
when 16#004C3# => romdata <= X"BA02001D";
when 16#004C4# => romdata <= X"85288001";
when 16#004C5# => romdata <= X"86006020";
when 16#004C6# => romdata <= X"88110002";
when 16#004C7# => romdata <= X"8728E002";
when 16#004C8# => romdata <= X"F4276088";
when 16#004C9# => romdata <= X"86020003";
when 16#004CA# => romdata <= X"C8222188";
when 16#004CB# => romdata <= X"80A72002";
when 16#004CC# => romdata <= X"02800009";
when 16#004CD# => romdata <= X"F620E088";
when 16#004CE# => romdata <= X"84006002";
when 16#004CF# => romdata <= X"82006001";
when 16#004D0# => romdata <= X"8528A002";
when 16#004D1# => romdata <= X"C2222004";
when 16#004D2# => romdata <= X"F2220002";
when 16#004D3# => romdata <= X"81C7E008";
when 16#004D4# => romdata <= X"91E82000";
when 16#004D5# => romdata <= X"C602218C";
when 16#004D6# => romdata <= X"8410C002";
when 16#004D7# => romdata <= X"10BFFFF7";
when 16#004D8# => romdata <= X"C422218C";
when 16#004D9# => romdata <= X"9007614C";
when 16#004DA# => romdata <= X"10BFFFCD";
when 16#004DB# => romdata <= X"D0276148";
when 16#004DC# => romdata <= X"81C3E008";
when 16#004DD# => romdata <= X"01000000";
when 16#004DE# => romdata <= X"81C3E008";
when 16#004DF# => romdata <= X"01000000";
when 16#004E0# => romdata <= X"81C3E008";
when 16#004E1# => romdata <= X"01000000";
when 16#004E2# => romdata <= X"82102001";
when 16#004E3# => romdata <= X"91D02000";
when 16#004E4# => romdata <= X"81C3E008";
when 16#004E5# => romdata <= X"01000000";
when 16#004E6# => romdata <= X"01000000";
when 16#004E7# => romdata <= X"A7580000";
when 16#004E8# => romdata <= X"A1480000";
when 16#004E9# => romdata <= X"A60CEFF0";
when 16#004EA# => romdata <= X"A734E004";
when 16#004EB# => romdata <= X"2B100008";
when 16#004EC# => romdata <= X"AA156280";
when 16#004ED# => romdata <= X"AC100013";
when 16#004EE# => romdata <= X"E8054000";
when 16#004EF# => romdata <= X"80A50016";
when 16#004F0# => romdata <= X"34800007";
when 16#004F1# => romdata <= X"AA05600C";
when 16#004F2# => romdata <= X"E6056004";
when 16#004F3# => romdata <= X"80A4C016";
when 16#004F4# => romdata <= X"36800013";
when 16#004F5# => romdata <= X"E6056008";
when 16#004F6# => romdata <= X"AA05600C";
when 16#004F7# => romdata <= X"E6054000";
when 16#004F8# => romdata <= X"A894E000";
when 16#004F9# => romdata <= X"12BFFFF7";
when 16#004FA# => romdata <= X"80A50016";
when 16#004FB# => romdata <= X"E6056004";
when 16#004FC# => romdata <= X"80A4E000";
when 16#004FD# => romdata <= X"12BFFFF3";
when 16#004FE# => romdata <= X"80A50016";
when 16#004FF# => romdata <= X"E6056008";
when 16#00500# => romdata <= X"80A4E000";
when 16#00501# => romdata <= X"12BFFFEF";
when 16#00502# => romdata <= X"80A50016";
when 16#00503# => romdata <= X"91D02000";
when 16#00504# => romdata <= X"01000000";
when 16#00505# => romdata <= X"01000000";
when 16#00506# => romdata <= X"01000000";
when 16#00507# => romdata <= X"81C4C000";
when 16#00508# => romdata <= X"01000000";
when 16#00509# => romdata <= X"01000000";
when 16#0050A# => romdata <= X"A7480000";
when 16#0050B# => romdata <= X"8B34E018";
when 16#0050C# => romdata <= X"8A096003";
when 16#0050D# => romdata <= X"80A16003";
when 16#0050E# => romdata <= X"12800011";
when 16#0050F# => romdata <= X"01000000";
when 16#00510# => romdata <= X"8B444000";
when 16#00511# => romdata <= X"03000008";
when 16#00512# => romdata <= X"8A114001";
when 16#00513# => romdata <= X"A3800005";
when 16#00514# => romdata <= X"01000000";
when 16#00515# => romdata <= X"01000000";
when 16#00516# => romdata <= X"01000000";
when 16#00517# => romdata <= X"8B444000";
when 16#00518# => romdata <= X"80894001";
when 16#00519# => romdata <= X"02800006";
when 16#0051A# => romdata <= X"01000000";
when 16#0051B# => romdata <= X"27100007";
when 16#0051C# => romdata <= X"A614E044";
when 16#0051D# => romdata <= X"81C4C000";
when 16#0051E# => romdata <= X"01000000";
when 16#0051F# => romdata <= X"91D02000";
when 16#00520# => romdata <= X"01000000";
when 16#00521# => romdata <= X"9DE3BFA0";
when 16#00522# => romdata <= X"3B100008";
when 16#00523# => romdata <= X"39100008";
when 16#00524# => romdata <= X"BA176270";
when 16#00525# => romdata <= X"B8172270";
when 16#00526# => romdata <= X"80A7401C";
when 16#00527# => romdata <= X"1A80000B";
when 16#00528# => romdata <= X"01000000";
when 16#00529# => romdata <= X"D0074000";
when 16#0052A# => romdata <= X"80A22000";
when 16#0052B# => romdata <= X"02800004";
when 16#0052C# => romdata <= X"BA076004";
when 16#0052D# => romdata <= X"9FC20000";
when 16#0052E# => romdata <= X"01000000";
when 16#0052F# => romdata <= X"80A7401C";
when 16#00530# => romdata <= X"2ABFFFFA";
when 16#00531# => romdata <= X"D0074000";
when 16#00532# => romdata <= X"81C7E008";
when 16#00533# => romdata <= X"81E80000";
when 16#00534# => romdata <= X"A7500000";
when 16#00535# => romdata <= X"AE100001";
when 16#00536# => romdata <= X"8334E001";
when 16#00537# => romdata <= X"2910000A";
when 16#00538# => romdata <= X"E805235C";
when 16#00539# => romdata <= X"A92CC014";
when 16#0053A# => romdata <= X"82150001";
when 16#0053B# => romdata <= X"81E00000";
when 16#0053C# => romdata <= X"81900001";
when 16#0053D# => romdata <= X"01000000";
when 16#0053E# => romdata <= X"01000000";
when 16#0053F# => romdata <= X"01000000";
when 16#00540# => romdata <= X"E03BA000";
when 16#00541# => romdata <= X"E43BA008";
when 16#00542# => romdata <= X"E83BA010";
when 16#00543# => romdata <= X"EC3BA018";
when 16#00544# => romdata <= X"F03BA020";
when 16#00545# => romdata <= X"F43BA028";
when 16#00546# => romdata <= X"F83BA030";
when 16#00547# => romdata <= X"FC3BA038";
when 16#00548# => romdata <= X"81E80000";
when 16#00549# => romdata <= X"82100017";
when 16#0054A# => romdata <= X"81C44000";
when 16#0054B# => romdata <= X"81CC8000";
when 16#0054C# => romdata <= X"01000000";
when 16#0054D# => romdata <= X"01000000";
when 16#0054E# => romdata <= X"01000000";
when 16#0054F# => romdata <= X"A7500000";
when 16#00550# => romdata <= X"A92CE001";
when 16#00551# => romdata <= X"2B10000A";
when 16#00552# => romdata <= X"EA05635C";
when 16#00553# => romdata <= X"AB34C015";
when 16#00554# => romdata <= X"AA154014";
when 16#00555# => romdata <= X"81900015";
when 16#00556# => romdata <= X"01000000";
when 16#00557# => romdata <= X"01000000";
when 16#00558# => romdata <= X"01000000";
when 16#00559# => romdata <= X"81E80000";
when 16#0055A# => romdata <= X"81E80000";
when 16#0055B# => romdata <= X"E01BA000";
when 16#0055C# => romdata <= X"E41BA008";
when 16#0055D# => romdata <= X"E81BA010";
when 16#0055E# => romdata <= X"EC1BA018";
when 16#0055F# => romdata <= X"F01BA020";
when 16#00560# => romdata <= X"F41BA028";
when 16#00561# => romdata <= X"F81BA030";
when 16#00562# => romdata <= X"FC1BA038";
when 16#00563# => romdata <= X"81E00000";
when 16#00564# => romdata <= X"81E00000";
when 16#00565# => romdata <= X"81C44000";
when 16#00566# => romdata <= X"81CC8000";
when 16#00567# => romdata <= X"A7500000";
when 16#00568# => romdata <= X"29100007";
when 16#00569# => romdata <= X"ADC52180";
when 16#0056A# => romdata <= X"01000000";
when 16#0056B# => romdata <= X"2710000A";
when 16#0056C# => romdata <= X"A614E294";
when 16#0056D# => romdata <= X"E024C000";
when 16#0056E# => romdata <= X"818C2020";
when 16#0056F# => romdata <= X"01000000";
when 16#00570# => romdata <= X"01000000";
when 16#00571# => romdata <= X"01000000";
when 16#00572# => romdata <= X"9DE3BFA0";
when 16#00573# => romdata <= X"9DE3BFA0";
when 16#00574# => romdata <= X"9DE3BFA0";
when 16#00575# => romdata <= X"9DE3BFA0";
when 16#00576# => romdata <= X"9DE3BFA0";
when 16#00577# => romdata <= X"9DE3BFA0";
when 16#00578# => romdata <= X"9DE3BFA0";
when 16#00579# => romdata <= X"81E80000";
when 16#0057A# => romdata <= X"81E80000";
when 16#0057B# => romdata <= X"81E80000";
when 16#0057C# => romdata <= X"81E80000";
when 16#0057D# => romdata <= X"81E80000";
when 16#0057E# => romdata <= X"81E80000";
when 16#0057F# => romdata <= X"81E80000";
when 16#00580# => romdata <= X"2710000A";
when 16#00581# => romdata <= X"A614E294";
when 16#00582# => romdata <= X"C024C000";
when 16#00583# => romdata <= X"E203A068";
when 16#00584# => romdata <= X"A4046004";
when 16#00585# => romdata <= X"E223A064";
when 16#00586# => romdata <= X"E423A068";
when 16#00587# => romdata <= X"10800204";
when 16#00588# => romdata <= X"AC100000";
when 16#00589# => romdata <= X"2910000A";
when 16#0058A# => romdata <= X"A8152278";
when 16#0058B# => romdata <= X"C2252000";
when 16#0058C# => romdata <= X"C8252004";
when 16#0058D# => romdata <= X"E0252010";
when 16#0058E# => romdata <= X"E2252014";
when 16#0058F# => romdata <= X"E4252018";
when 16#00590# => romdata <= X"E825201C";
when 16#00591# => romdata <= X"81E80000";
when 16#00592# => romdata <= X"83480000";
when 16#00593# => romdata <= X"82106F00";
when 16#00594# => romdata <= X"81886020";
when 16#00595# => romdata <= X"01000000";
when 16#00596# => romdata <= X"01000000";
when 16#00597# => romdata <= X"01000000";
when 16#00598# => romdata <= X"0910000A";
when 16#00599# => romdata <= X"C801235C";
when 16#0059A# => romdata <= X"81E00000";
when 16#0059B# => romdata <= X"88212001";
when 16#0059C# => romdata <= X"80A920FF";
when 16#0059D# => romdata <= X"02800003";
when 16#0059E# => romdata <= X"01000000";
when 16#0059F# => romdata <= X"01000000";
when 16#005A0# => romdata <= X"80A10000";
when 16#005A1# => romdata <= X"12BFFFF9";
when 16#005A2# => romdata <= X"01000000";
when 16#005A3# => romdata <= X"0910000A";
when 16#005A4# => romdata <= X"C801235C";
when 16#005A5# => romdata <= X"81E80000";
when 16#005A6# => romdata <= X"80A920FF";
when 16#005A7# => romdata <= X"02800003";
when 16#005A8# => romdata <= X"01000000";
when 16#005A9# => romdata <= X"01000000";
when 16#005AA# => romdata <= X"88212001";
when 16#005AB# => romdata <= X"80A10000";
when 16#005AC# => romdata <= X"12BFFFF9";
when 16#005AD# => romdata <= X"01000000";
when 16#005AE# => romdata <= X"81E00000";
when 16#005AF# => romdata <= X"2910000A";
when 16#005B0# => romdata <= X"A8152278";
when 16#005B1# => romdata <= X"C8052004";
when 16#005B2# => romdata <= X"C2052000";
when 16#005B3# => romdata <= X"E0052010";
when 16#005B4# => romdata <= X"E2052014";
when 16#005B5# => romdata <= X"E4052018";
when 16#005B6# => romdata <= X"C025201C";
when 16#005B7# => romdata <= X"818C2000";
when 16#005B8# => romdata <= X"01000000";
when 16#005B9# => romdata <= X"01000000";
when 16#005BA# => romdata <= X"01000000";
when 16#005BB# => romdata <= X"81C48000";
when 16#005BC# => romdata <= X"81CCA004";
when 16#005BD# => romdata <= X"A0142F00";
when 16#005BE# => romdata <= X"81880010";
when 16#005BF# => romdata <= X"01000000";
when 16#005C0# => romdata <= X"01000000";
when 16#005C1# => romdata <= X"01000000";
when 16#005C2# => romdata <= X"81C48000";
when 16#005C3# => romdata <= X"81CCA004";
when 16#005C4# => romdata <= X"80A66002";
when 16#005C5# => romdata <= X"12800005";
when 16#005C6# => romdata <= X"A8142F00";
when 16#005C7# => romdata <= X"81880014";
when 16#005C8# => romdata <= X"B0142020";
when 16#005C9# => romdata <= X"3080001F";
when 16#005CA# => romdata <= X"80A66003";
when 16#005CB# => romdata <= X"12800006";
when 16#005CC# => romdata <= X"A80E2F00";
when 16#005CD# => romdata <= X"AA2C2F00";
when 16#005CE# => romdata <= X"A8154014";
when 16#005CF# => romdata <= X"81880014";
when 16#005D0# => romdata <= X"30800018";
when 16#005D1# => romdata <= X"80A66004";
when 16#005D2# => romdata <= X"12800008";
when 16#005D3# => romdata <= X"A9480000";
when 16#005D4# => romdata <= X"A8152040";
when 16#005D5# => romdata <= X"81880014";
when 16#005D6# => romdata <= X"01000000";
when 16#005D7# => romdata <= X"01000000";
when 16#005D8# => romdata <= X"01000000";
when 16#005D9# => romdata <= X"3080000F";
when 16#005DA# => romdata <= X"80A66005";
when 16#005DB# => romdata <= X"12800008";
when 16#005DC# => romdata <= X"A9480000";
when 16#005DD# => romdata <= X"A82D2040";
when 16#005DE# => romdata <= X"81880014";
when 16#005DF# => romdata <= X"01000000";
when 16#005E0# => romdata <= X"01000000";
when 16#005E1# => romdata <= X"01000000";
when 16#005E2# => romdata <= X"30800006";
when 16#005E3# => romdata <= X"80A66006";
when 16#005E4# => romdata <= X"12800003";
when 16#005E5# => romdata <= X"01000000";
when 16#005E6# => romdata <= X"30BFFFA3";
when 16#005E7# => romdata <= X"91D02000";
when 16#005E8# => romdata <= X"81C48000";
when 16#005E9# => romdata <= X"81CCA004";
when 16#005EA# => romdata <= X"92102003";
when 16#005EB# => romdata <= X"81C3E008";
when 16#005EC# => romdata <= X"91D02002";
when 16#005ED# => romdata <= X"92102002";
when 16#005EE# => romdata <= X"81C3E008";
when 16#005EF# => romdata <= X"91D02002";
when 16#005F0# => romdata <= X"92102006";
when 16#005F1# => romdata <= X"81C3E008";
when 16#005F2# => romdata <= X"91D02002";
when 16#005F3# => romdata <= X"27000004";
when 16#005F4# => romdata <= X"A0140013";
when 16#005F5# => romdata <= X"A6142F00";
when 16#005F6# => romdata <= X"818CE000";
when 16#005F7# => romdata <= X"01000000";
when 16#005F8# => romdata <= X"01000000";
when 16#005F9# => romdata <= X"01000000";
when 16#005FA# => romdata <= X"A7480000";
when 16#005FB# => romdata <= X"29000004";
when 16#005FC# => romdata <= X"A68CC014";
when 16#005FD# => romdata <= X"12800003";
when 16#005FE# => romdata <= X"01000000";
when 16#005FF# => romdata <= X"91D02000";
when 16#00600# => romdata <= X"2910000A";
when 16#00601# => romdata <= X"A815233C";
when 16#00602# => romdata <= X"E8050000";
when 16#00603# => romdata <= X"2B10000A";
when 16#00604# => romdata <= X"AA156338";
when 16#00605# => romdata <= X"EA054000";
when 16#00606# => romdata <= X"80A50015";
when 16#00607# => romdata <= X"0280002D";
when 16#00608# => romdata <= X"01000000";
when 16#00609# => romdata <= X"80A00015";
when 16#0060A# => romdata <= X"02800013";
when 16#0060B# => romdata <= X"01000000";
when 16#0060C# => romdata <= X"C13D6000";
when 16#0060D# => romdata <= X"C53D6008";
when 16#0060E# => romdata <= X"C93D6010";
when 16#0060F# => romdata <= X"CD3D6018";
when 16#00610# => romdata <= X"D13D6020";
when 16#00611# => romdata <= X"D53D6028";
when 16#00612# => romdata <= X"D93D6030";
when 16#00613# => romdata <= X"DD3D6038";
when 16#00614# => romdata <= X"E13D6040";
when 16#00615# => romdata <= X"E53D6048";
when 16#00616# => romdata <= X"E93D6050";
when 16#00617# => romdata <= X"ED3D6058";
when 16#00618# => romdata <= X"F13D6060";
when 16#00619# => romdata <= X"F53D6068";
when 16#0061A# => romdata <= X"F93D6070";
when 16#0061B# => romdata <= X"FD3D6078";
when 16#0061C# => romdata <= X"C12D6080";
when 16#0061D# => romdata <= X"2D10000A";
when 16#0061E# => romdata <= X"AC15A338";
when 16#0061F# => romdata <= X"E8258000";
when 16#00620# => romdata <= X"80A00014";
when 16#00621# => romdata <= X"02800013";
when 16#00622# => romdata <= X"01000000";
when 16#00623# => romdata <= X"C11D2000";
when 16#00624# => romdata <= X"C51D2008";
when 16#00625# => romdata <= X"C91D2010";
when 16#00626# => romdata <= X"CD1D2018";
when 16#00627# => romdata <= X"D11D2020";
when 16#00628# => romdata <= X"D51D2028";
when 16#00629# => romdata <= X"D91D2030";
when 16#0062A# => romdata <= X"DD1D2038";
when 16#0062B# => romdata <= X"E11D2040";
when 16#0062C# => romdata <= X"E51D2048";
when 16#0062D# => romdata <= X"E91D2050";
when 16#0062E# => romdata <= X"ED1D2058";
when 16#0062F# => romdata <= X"F11D2060";
when 16#00630# => romdata <= X"F51D2068";
when 16#00631# => romdata <= X"F91D2070";
when 16#00632# => romdata <= X"FD1D2078";
when 16#00633# => romdata <= X"C10D2080";
when 16#00634# => romdata <= X"818C2000";
when 16#00635# => romdata <= X"01000000";
when 16#00636# => romdata <= X"01000000";
when 16#00637# => romdata <= X"01000000";
when 16#00638# => romdata <= X"81C44000";
when 16#00639# => romdata <= X"81CC8000";
when 16#0063A# => romdata <= X"AE25A010";
when 16#0063B# => romdata <= X"A7500000";
when 16#0063C# => romdata <= X"2D100006";
when 16#0063D# => romdata <= X"AC15A0FC";
when 16#0063E# => romdata <= X"29100007";
when 16#0063F# => romdata <= X"81C52348";
when 16#00640# => romdata <= X"01000000";
when 16#00641# => romdata <= X"1110000A";
when 16#00642# => romdata <= X"90122348";
when 16#00643# => romdata <= X"D2020000";
when 16#00644# => romdata <= X"92026001";
when 16#00645# => romdata <= X"D2220000";
when 16#00646# => romdata <= X"932DE008";
when 16#00647# => romdata <= X"902C2F00";
when 16#00648# => romdata <= X"92120009";
when 16#00649# => romdata <= X"1110000A";
when 16#0064A# => romdata <= X"90122340";
when 16#0064B# => romdata <= X"D0020000";
when 16#0064C# => romdata <= X"80A00008";
when 16#0064D# => romdata <= X"22800002";
when 16#0064E# => romdata <= X"92126F00";
when 16#0064F# => romdata <= X"818A6020";
when 16#00650# => romdata <= X"01000000";
when 16#00651# => romdata <= X"01000000";
when 16#00652# => romdata <= X"01000000";
when 16#00653# => romdata <= X"90100017";
when 16#00654# => romdata <= X"40000037";
when 16#00655# => romdata <= X"9203A0F8";
when 16#00656# => romdata <= X"92142F00";
when 16#00657# => romdata <= X"818A6020";
when 16#00658# => romdata <= X"01000000";
when 16#00659# => romdata <= X"01000000";
when 16#0065A# => romdata <= X"01000000";
when 16#0065B# => romdata <= X"1110000A";
when 16#0065C# => romdata <= X"90122348";
when 16#0065D# => romdata <= X"D2020000";
when 16#0065E# => romdata <= X"92226001";
when 16#0065F# => romdata <= X"D2220000";
when 16#00660# => romdata <= X"1080019A";
when 16#00661# => romdata <= X"AC100000";
when 16#00662# => romdata <= X"9DE3BFA0";
when 16#00663# => romdata <= X"0510000B";
when 16#00664# => romdata <= X"832E6002";
when 16#00665# => romdata <= X"8410A238";
when 16#00666# => romdata <= X"88102000";
when 16#00667# => romdata <= X"80A6601F";
when 16#00668# => romdata <= X"14800017";
when 16#00669# => romdata <= X"DE008001";
when 16#0066A# => romdata <= X"B32E6004";
when 16#0066B# => romdata <= X"1B10000B";
when 16#0066C# => romdata <= X"80A3E000";
when 16#0066D# => romdata <= X"9A136038";
when 16#0066E# => romdata <= X"0280000D";
when 16#0066F# => romdata <= X"8806400D";
when 16#00670# => romdata <= X"80A3C004";
when 16#00671# => romdata <= X"12800006";
when 16#00672# => romdata <= X"8610000F";
when 16#00673# => romdata <= X"1080000E";
when 16#00674# => romdata <= X"C800C000";
when 16#00675# => romdata <= X"2280000C";
when 16#00676# => romdata <= X"C800C000";
when 16#00677# => romdata <= X"C600E00C";
when 16#00678# => romdata <= X"80A0E000";
when 16#00679# => romdata <= X"12BFFFFC";
when 16#0067A# => romdata <= X"80A10003";
when 16#0067B# => romdata <= X"F026400D";
when 16#0067C# => romdata <= X"DE21200C";
when 16#0067D# => romdata <= X"C8208001";
when 16#0067E# => romdata <= X"88102000";
when 16#0067F# => romdata <= X"81C7E008";
when 16#00680# => romdata <= X"91E80004";
when 16#00681# => romdata <= X"F020C000";
when 16#00682# => romdata <= X"81C7E008";
when 16#00683# => romdata <= X"91E80004";
when 16#00684# => romdata <= X"912A2002";
when 16#00685# => romdata <= X"0310000B";
when 16#00686# => romdata <= X"82106238";
when 16#00687# => romdata <= X"C4004008";
when 16#00688# => romdata <= X"C422600C";
when 16#00689# => romdata <= X"81C3E008";
when 16#0068A# => romdata <= X"D2204008";
when 16#0068B# => romdata <= X"9DE3BFA0";
when 16#0068C# => romdata <= X"0510000A";
when 16#0068D# => romdata <= X"8210A34C";
when 16#0068E# => romdata <= X"C2006004";
when 16#0068F# => romdata <= X"80A04018";
when 16#00690# => romdata <= X"22800039";
when 16#00691# => romdata <= X"C400A34C";
when 16#00692# => romdata <= X"80A62000";
when 16#00693# => romdata <= X"22800002";
when 16#00694# => romdata <= X"B0100001";
when 16#00695# => romdata <= X"B72E2002";
when 16#00696# => romdata <= X"0310000B";
when 16#00697# => romdata <= X"82106238";
when 16#00698# => romdata <= X"FA00401B";
when 16#00699# => romdata <= X"80A76000";
when 16#0069A# => romdata <= X"0280002D";
when 16#0069B# => romdata <= X"3510000B";
when 16#0069C# => romdata <= X"2510000A";
when 16#0069D# => romdata <= X"2310000A";
when 16#0069E# => romdata <= X"1080001C";
when 16#0069F# => romdata <= X"2110000A";
when 16#006A0# => romdata <= X"C607001B";
when 16#006A1# => romdata <= X"8600E001";
when 16#006A2# => romdata <= X"C404A3B0";
when 16#006A3# => romdata <= X"80A0A000";
when 16#006A4# => romdata <= X"02800005";
when 16#006A5# => romdata <= X"C627001B";
when 16#006A6# => romdata <= X"9FC08000";
when 16#006A7# => romdata <= X"01000000";
when 16#006A8# => romdata <= X"C2074000";
when 16#006A9# => romdata <= X"D2076008";
when 16#006AA# => romdata <= X"90100018";
when 16#006AB# => romdata <= X"9FC04000";
when 16#006AC# => romdata <= X"94100019";
when 16#006AD# => romdata <= X"C20463AC";
when 16#006AE# => romdata <= X"80A06000";
when 16#006AF# => romdata <= X"22800005";
when 16#006B0# => romdata <= X"C207001B";
when 16#006B1# => romdata <= X"9FC04000";
when 16#006B2# => romdata <= X"01000000";
when 16#006B3# => romdata <= X"C207001B";
when 16#006B4# => romdata <= X"82007FFF";
when 16#006B5# => romdata <= X"C227001B";
when 16#006B6# => romdata <= X"FA07600C";
when 16#006B7# => romdata <= X"80A76000";
when 16#006B8# => romdata <= X"0280000F";
when 16#006B9# => romdata <= X"01000000";
when 16#006BA# => romdata <= X"C2074000";
when 16#006BB# => romdata <= X"80A06000";
when 16#006BC# => romdata <= X"02BFFFFA";
when 16#006BD# => romdata <= X"C406A034";
when 16#006BE# => romdata <= X"80A0A000";
when 16#006BF# => romdata <= X"12BFFFE1";
when 16#006C0# => romdata <= X"B81423B4";
when 16#006C1# => romdata <= X"C407001B";
when 16#006C2# => romdata <= X"80A0A000";
when 16#006C3# => romdata <= X"32BFFFF4";
when 16#006C4# => romdata <= X"FA07600C";
when 16#006C5# => romdata <= X"10BFFFDC";
when 16#006C6# => romdata <= X"86102000";
when 16#006C7# => romdata <= X"81C7E008";
when 16#006C8# => romdata <= X"81E80000";
when 16#006C9# => romdata <= X"F000A0C0";
when 16#006CA# => romdata <= X"10BFFFC8";
when 16#006CB# => romdata <= X"B00E201F";
when 16#006CC# => romdata <= X"8C10000F";
when 16#006CD# => romdata <= X"A7480000";
when 16#006CE# => romdata <= X"8B34E018";
when 16#006CF# => romdata <= X"8A09600F";
when 16#006D0# => romdata <= X"80A16003";
when 16#006D1# => romdata <= X"02800002";
when 16#006D2# => romdata <= X"10800039";
when 16#006D3# => romdata <= X"90102001";
when 16#006D4# => romdata <= X"92102006";
when 16#006D5# => romdata <= X"4000016E";
when 16#006D6# => romdata <= X"01000000";
when 16#006D7# => romdata <= X"80A00008";
when 16#006D8# => romdata <= X"02800033";
when 16#006D9# => romdata <= X"01000000";
when 16#006DA# => romdata <= X"C2022010";
when 16#006DB# => romdata <= X"113FFC00";
when 16#006DC# => romdata <= X"82084008";
when 16#006DD# => romdata <= X"110003FC";
when 16#006DE# => romdata <= X"84104008";
when 16#006DF# => romdata <= X"90100002";
when 16#006E0# => romdata <= X"92102001";
when 16#006E1# => romdata <= X"9410200C";
when 16#006E2# => romdata <= X"40000177";
when 16#006E3# => romdata <= X"01000000";
when 16#006E4# => romdata <= X"80A00008";
when 16#006E5# => romdata <= X"02800026";
when 16#006E6# => romdata <= X"01000000";
when 16#006E7# => romdata <= X"40000187";
when 16#006E8# => romdata <= X"92100001";
when 16#006E9# => romdata <= X"0B10000A";
when 16#006EA# => romdata <= X"8A116354";
when 16#006EB# => romdata <= X"D2214000";
when 16#006EC# => romdata <= X"90100002";
when 16#006ED# => romdata <= X"92102001";
when 16#006EE# => romdata <= X"94102011";
when 16#006EF# => romdata <= X"4000016A";
when 16#006F0# => romdata <= X"01000000";
when 16#006F1# => romdata <= X"80A00008";
when 16#006F2# => romdata <= X"02800019";
when 16#006F3# => romdata <= X"01000000";
when 16#006F4# => romdata <= X"4000017A";
when 16#006F5# => romdata <= X"92100001";
when 16#006F6# => romdata <= X"92026010";
when 16#006F7# => romdata <= X"0B10000A";
when 16#006F8# => romdata <= X"8A116370";
when 16#006F9# => romdata <= X"D2214000";
when 16#006FA# => romdata <= X"90100002";
when 16#006FB# => romdata <= X"92102001";
when 16#006FC# => romdata <= X"9410200D";
when 16#006FD# => romdata <= X"4000015C";
when 16#006FE# => romdata <= X"01000000";
when 16#006FF# => romdata <= X"80A00008";
when 16#00700# => romdata <= X"0280000B";
when 16#00701# => romdata <= X"01000000";
when 16#00702# => romdata <= X"4000016C";
when 16#00703# => romdata <= X"92100001";
when 16#00704# => romdata <= X"0B10000A";
when 16#00705# => romdata <= X"8A11634C";
when 16#00706# => romdata <= X"D2214000";
when 16#00707# => romdata <= X"D4026010";
when 16#00708# => romdata <= X"9532A010";
when 16#00709# => romdata <= X"940AA00F";
when 16#0070A# => romdata <= X"D4216004";
when 16#0070B# => romdata <= X"9E100006";
when 16#0070C# => romdata <= X"81C3E008";
when 16#0070D# => romdata <= X"01000000";
when 16#0070E# => romdata <= X"0310000A";
when 16#0070F# => romdata <= X"82106368";
when 16#00710# => romdata <= X"01000000";
when 16#00711# => romdata <= X"03100007";
when 16#00712# => romdata <= X"821060F8";
when 16#00713# => romdata <= X"9FC04000";
when 16#00714# => romdata <= X"01000000";
when 16#00715# => romdata <= X"03100000";
when 16#00716# => romdata <= X"82106000";
when 16#00717# => romdata <= X"81980001";
when 16#00718# => romdata <= X"03100007";
when 16#00719# => romdata <= X"82106160";
when 16#0071A# => romdata <= X"9FC04000";
when 16#0071B# => romdata <= X"01000000";
when 16#0071C# => romdata <= X"03100007";
when 16#0071D# => romdata <= X"821060E8";
when 16#0071E# => romdata <= X"9FC04000";
when 16#0071F# => romdata <= X"01000000";
when 16#00720# => romdata <= X"8B444000";
when 16#00721# => romdata <= X"8B31601C";
when 16#00722# => romdata <= X"80A14000";
when 16#00723# => romdata <= X"12800006";
when 16#00724# => romdata <= X"01000000";
when 16#00725# => romdata <= X"7FFFFFA7";
when 16#00726# => romdata <= X"01000000";
when 16#00727# => romdata <= X"7FFFF942";
when 16#00728# => romdata <= X"01000000";
when 16#00729# => romdata <= X"9C23A040";
when 16#0072A# => romdata <= X"7FFFF8D9";
when 16#0072B# => romdata <= X"01000000";
when 16#0072C# => romdata <= X"82102001";
when 16#0072D# => romdata <= X"91D02000";
when 16#0072E# => romdata <= X"01000000";
when 16#0072F# => romdata <= X"29000004";
when 16#00730# => romdata <= X"A68C0014";
when 16#00731# => romdata <= X"32800003";
when 16#00732# => romdata <= X"A02C0014";
when 16#00733# => romdata <= X"91D02000";
when 16#00734# => romdata <= X"81880010";
when 16#00735# => romdata <= X"01000000";
when 16#00736# => romdata <= X"01000000";
when 16#00737# => romdata <= X"01000000";
when 16#00738# => romdata <= X"81C48000";
when 16#00739# => romdata <= X"81CCA004";
when 16#0073A# => romdata <= X"81C3E008";
when 16#0073B# => romdata <= X"01000000";
when 16#0073C# => romdata <= X"81C1E008";
when 16#0073D# => romdata <= X"01000000";
when 16#0073E# => romdata <= X"A7480000";
when 16#0073F# => romdata <= X"8B34E018";
when 16#00740# => romdata <= X"8A096003";
when 16#00741# => romdata <= X"80A16003";
when 16#00742# => romdata <= X"12800008";
when 16#00743# => romdata <= X"01000000";
when 16#00744# => romdata <= X"2110000A";
when 16#00745# => romdata <= X"A0142364";
when 16#00746# => romdata <= X"A2102003";
when 16#00747# => romdata <= X"E2240000";
when 16#00748# => romdata <= X"8B444000";
when 16#00749# => romdata <= X"10800001";
when 16#0074A# => romdata <= X"8A09601F";
when 16#0074B# => romdata <= X"2710000A";
when 16#0074C# => romdata <= X"A614E35C";
when 16#0074D# => romdata <= X"CA24C000";
when 16#0074E# => romdata <= X"8A016001";
when 16#0074F# => romdata <= X"2710000A";
when 16#00750# => romdata <= X"A614E358";
when 16#00751# => romdata <= X"CA24C000";
when 16#00752# => romdata <= X"2710000A";
when 16#00753# => romdata <= X"A614E360";
when 16#00754# => romdata <= X"8A216002";
when 16#00755# => romdata <= X"CA24C000";
when 16#00756# => romdata <= X"81C3E008";
when 16#00757# => romdata <= X"01000000";
when 16#00758# => romdata <= X"81C3E008";
when 16#00759# => romdata <= X"01000000";
when 16#0075A# => romdata <= X"91D02000";
when 16#0075B# => romdata <= X"01000000";
when 16#0075C# => romdata <= X"01000000";
when 16#0075D# => romdata <= X"01000000";
when 16#0075E# => romdata <= X"81C44000";
when 16#0075F# => romdata <= X"81CC8000";
when 16#00760# => romdata <= X"AA27A140";
when 16#00761# => romdata <= X"E0256060";
when 16#00762# => romdata <= X"E2256064";
when 16#00763# => romdata <= X"E4256068";
when 16#00764# => romdata <= X"C2256074";
when 16#00765# => romdata <= X"C43D6078";
when 16#00766# => romdata <= X"C83D6080";
when 16#00767# => romdata <= X"CC3D6088";
when 16#00768# => romdata <= X"85400000";
when 16#00769# => romdata <= X"C425606C";
when 16#0076A# => romdata <= X"F03D6090";
when 16#0076B# => romdata <= X"F43D6098";
when 16#0076C# => romdata <= X"F83D60A0";
when 16#0076D# => romdata <= X"FC3D60A8";
when 16#0076E# => romdata <= X"0510000A";
when 16#0076F# => romdata <= X"C600A33C";
when 16#00770# => romdata <= X"C625613C";
when 16#00771# => romdata <= X"860560B0";
when 16#00772# => romdata <= X"C620A33C";
when 16#00773# => romdata <= X"A8102001";
when 16#00774# => romdata <= X"A92D0010";
when 16#00775# => romdata <= X"808D0013";
when 16#00776# => romdata <= X"02800013";
when 16#00777# => romdata <= X"01000000";
when 16#00778# => romdata <= X"8534E001";
when 16#00779# => romdata <= X"0710000A";
when 16#0077A# => romdata <= X"C600E35C";
when 16#0077B# => romdata <= X"A72CC003";
when 16#0077C# => romdata <= X"8414C002";
when 16#0077D# => romdata <= X"8408A0FF";
when 16#0077E# => romdata <= X"81E00000";
when 16#0077F# => romdata <= X"8190A000";
when 16#00780# => romdata <= X"E03BA000";
when 16#00781# => romdata <= X"E43BA008";
when 16#00782# => romdata <= X"E83BA010";
when 16#00783# => romdata <= X"EC3BA018";
when 16#00784# => romdata <= X"F03BA020";
when 16#00785# => romdata <= X"F43BA028";
when 16#00786# => romdata <= X"F83BA030";
when 16#00787# => romdata <= X"FC3BA038";
when 16#00788# => romdata <= X"81E80000";
when 16#00789# => romdata <= X"81C5A008";
when 16#0078A# => romdata <= X"9C100015";
when 16#0078B# => romdata <= X"0510000A";
when 16#0078C# => romdata <= X"8410A3A8";
when 16#0078D# => romdata <= X"C4008000";
when 16#0078E# => romdata <= X"80A08000";
when 16#0078F# => romdata <= X"02800004";
when 16#00790# => romdata <= X"01000000";
when 16#00791# => romdata <= X"9FC08000";
when 16#00792# => romdata <= X"9203A0F8";
when 16#00793# => romdata <= X"C403A13C";
when 16#00794# => romdata <= X"0710000A";
when 16#00795# => romdata <= X"C420E33C";
when 16#00796# => romdata <= X"818C2000";
when 16#00797# => romdata <= X"82102002";
when 16#00798# => romdata <= X"83284010";
when 16#00799# => romdata <= X"0510000A";
when 16#0079A# => romdata <= X"C400A358";
when 16#0079B# => romdata <= X"85304002";
when 16#0079C# => romdata <= X"82104002";
when 16#0079D# => romdata <= X"85500000";
when 16#0079E# => romdata <= X"80888001";
when 16#0079F# => romdata <= X"02800020";
when 16#007A0# => romdata <= X"8328A001";
when 16#007A1# => romdata <= X"0710000A";
when 16#007A2# => romdata <= X"C600E35C";
when 16#007A3# => romdata <= X"85308003";
when 16#007A4# => romdata <= X"82104002";
when 16#007A5# => romdata <= X"820860FF";
when 16#007A6# => romdata <= X"81906000";
when 16#007A7# => romdata <= X"C203A06C";
when 16#007A8# => romdata <= X"81806000";
when 16#007A9# => romdata <= X"F01BA090";
when 16#007AA# => romdata <= X"F41BA098";
when 16#007AB# => romdata <= X"F81BA0A0";
when 16#007AC# => romdata <= X"FC1BA0A8";
when 16#007AD# => romdata <= X"C203A074";
when 16#007AE# => romdata <= X"C41BA078";
when 16#007AF# => romdata <= X"C81BA080";
when 16#007B0# => romdata <= X"CC1BA088";
when 16#007B1# => romdata <= X"E003A060";
when 16#007B2# => romdata <= X"E203A064";
when 16#007B3# => romdata <= X"E403A068";
when 16#007B4# => romdata <= X"81E80000";
when 16#007B5# => romdata <= X"E01BA000";
when 16#007B6# => romdata <= X"E41BA008";
when 16#007B7# => romdata <= X"E81BA010";
when 16#007B8# => romdata <= X"EC1BA018";
when 16#007B9# => romdata <= X"F01BA020";
when 16#007BA# => romdata <= X"F41BA028";
when 16#007BB# => romdata <= X"F81BA030";
when 16#007BC# => romdata <= X"FC1BA038";
when 16#007BD# => romdata <= X"1080000F";
when 16#007BE# => romdata <= X"81E00000";
when 16#007BF# => romdata <= X"C203A06C";
when 16#007C0# => romdata <= X"81806000";
when 16#007C1# => romdata <= X"F01BA090";
when 16#007C2# => romdata <= X"F41BA098";
when 16#007C3# => romdata <= X"F81BA0A0";
when 16#007C4# => romdata <= X"FC1BA0A8";
when 16#007C5# => romdata <= X"C203A074";
when 16#007C6# => romdata <= X"C41BA078";
when 16#007C7# => romdata <= X"C81BA080";
when 16#007C8# => romdata <= X"CC1BA088";
when 16#007C9# => romdata <= X"E003A060";
when 16#007CA# => romdata <= X"E203A064";
when 16#007CB# => romdata <= X"E403A068";
when 16#007CC# => romdata <= X"818C2000";
when 16#007CD# => romdata <= X"01000000";
when 16#007CE# => romdata <= X"01000000";
when 16#007CF# => romdata <= X"01000000";
when 16#007D0# => romdata <= X"81C44000";
when 16#007D1# => romdata <= X"81CC8000";
when 16#007D2# => romdata <= X"AA27A140";
when 16#007D3# => romdata <= X"E0256138";
when 16#007D4# => romdata <= X"29000004";
when 16#007D5# => romdata <= X"A02C0014";
when 16#007D6# => romdata <= X"C2256074";
when 16#007D7# => romdata <= X"C43D6078";
when 16#007D8# => romdata <= X"C83D6080";
when 16#007D9# => romdata <= X"CC3D6088";
when 16#007DA# => romdata <= X"85400000";
when 16#007DB# => romdata <= X"C425606C";
when 16#007DC# => romdata <= X"0510000A";
when 16#007DD# => romdata <= X"C600A33C";
when 16#007DE# => romdata <= X"C625613C";
when 16#007DF# => romdata <= X"860560B0";
when 16#007E0# => romdata <= X"C620A33C";
when 16#007E1# => romdata <= X"C020E080";
when 16#007E2# => romdata <= X"A8102001";
when 16#007E3# => romdata <= X"A92D0010";
when 16#007E4# => romdata <= X"808D0013";
when 16#007E5# => romdata <= X"02800013";
when 16#007E6# => romdata <= X"01000000";
when 16#007E7# => romdata <= X"8534E001";
when 16#007E8# => romdata <= X"0710000A";
when 16#007E9# => romdata <= X"C600E35C";
when 16#007EA# => romdata <= X"A72CC003";
when 16#007EB# => romdata <= X"8414C002";
when 16#007EC# => romdata <= X"8408A0FF";
when 16#007ED# => romdata <= X"81E00000";
when 16#007EE# => romdata <= X"8190A000";
when 16#007EF# => romdata <= X"E03BA000";
when 16#007F0# => romdata <= X"E43BA008";
when 16#007F1# => romdata <= X"E83BA010";
when 16#007F2# => romdata <= X"EC3BA018";
when 16#007F3# => romdata <= X"F03BA020";
when 16#007F4# => romdata <= X"F43BA028";
when 16#007F5# => romdata <= X"F83BA030";
when 16#007F6# => romdata <= X"FC3BA038";
when 16#007F7# => romdata <= X"81E80000";
when 16#007F8# => romdata <= X"81C5A008";
when 16#007F9# => romdata <= X"9C100015";
when 16#007FA# => romdata <= X"0510000A";
when 16#007FB# => romdata <= X"8410A3A8";
when 16#007FC# => romdata <= X"C4008000";
when 16#007FD# => romdata <= X"80A08000";
when 16#007FE# => romdata <= X"02800004";
when 16#007FF# => romdata <= X"01000000";
when 16#00800# => romdata <= X"9FC08000";
when 16#00801# => romdata <= X"9203A0F8";
when 16#00802# => romdata <= X"C403A13C";
when 16#00803# => romdata <= X"0710000A";
when 16#00804# => romdata <= X"C420E33C";
when 16#00805# => romdata <= X"0710000A";
when 16#00806# => romdata <= X"C600E338";
when 16#00807# => romdata <= X"80A08003";
when 16#00808# => romdata <= X"12800008";
when 16#00809# => romdata <= X"01000000";
when 16#0080A# => romdata <= X"C403A138";
when 16#0080B# => romdata <= X"07000004";
when 16#0080C# => romdata <= X"84088003";
when 16#0080D# => romdata <= X"A02C0003";
when 16#0080E# => romdata <= X"A0140002";
when 16#0080F# => romdata <= X"30800006";
when 16#00810# => romdata <= X"8403A0B0";
when 16#00811# => romdata <= X"80A08003";
when 16#00812# => romdata <= X"12800003";
when 16#00813# => romdata <= X"0710000A";
when 16#00814# => romdata <= X"C020E338";
when 16#00815# => romdata <= X"818C2000";
when 16#00816# => romdata <= X"82102002";
when 16#00817# => romdata <= X"83284010";
when 16#00818# => romdata <= X"0510000A";
when 16#00819# => romdata <= X"C400A358";
when 16#0081A# => romdata <= X"85304002";
when 16#0081B# => romdata <= X"82104002";
when 16#0081C# => romdata <= X"85500000";
when 16#0081D# => romdata <= X"80888001";
when 16#0081E# => romdata <= X"02800019";
when 16#0081F# => romdata <= X"8328A001";
when 16#00820# => romdata <= X"0710000A";
when 16#00821# => romdata <= X"C600E35C";
when 16#00822# => romdata <= X"85308003";
when 16#00823# => romdata <= X"82104002";
when 16#00824# => romdata <= X"820860FF";
when 16#00825# => romdata <= X"81906000";
when 16#00826# => romdata <= X"C203A06C";
when 16#00827# => romdata <= X"81806000";
when 16#00828# => romdata <= X"C203A074";
when 16#00829# => romdata <= X"C41BA078";
when 16#0082A# => romdata <= X"C81BA080";
when 16#0082B# => romdata <= X"CC1BA088";
when 16#0082C# => romdata <= X"81E80000";
when 16#0082D# => romdata <= X"E01BA000";
when 16#0082E# => romdata <= X"E41BA008";
when 16#0082F# => romdata <= X"E81BA010";
when 16#00830# => romdata <= X"EC1BA018";
when 16#00831# => romdata <= X"F01BA020";
when 16#00832# => romdata <= X"F41BA028";
when 16#00833# => romdata <= X"F81BA030";
when 16#00834# => romdata <= X"FC1BA038";
when 16#00835# => romdata <= X"10800008";
when 16#00836# => romdata <= X"81E00000";
when 16#00837# => romdata <= X"C203A06C";
when 16#00838# => romdata <= X"81806000";
when 16#00839# => romdata <= X"C203A074";
when 16#0083A# => romdata <= X"C41BA078";
when 16#0083B# => romdata <= X"C81BA080";
when 16#0083C# => romdata <= X"CC1BA088";
when 16#0083D# => romdata <= X"818C2000";
when 16#0083E# => romdata <= X"01000000";
when 16#0083F# => romdata <= X"01000000";
when 16#00840# => romdata <= X"01000000";
when 16#00841# => romdata <= X"81C44000";
when 16#00842# => romdata <= X"81CC8000";
when 16#00843# => romdata <= X"82100008";
when 16#00844# => romdata <= X"9A103800";
when 16#00845# => romdata <= X"96102000";
when 16#00846# => romdata <= X"912AE005";
when 16#00847# => romdata <= X"98034008";
when 16#00848# => romdata <= X"D4034008";
when 16#00849# => romdata <= X"9132A018";
when 16#0084A# => romdata <= X"80A20001";
when 16#0084B# => romdata <= X"32800008";
when 16#0084C# => romdata <= X"9602E001";
when 16#0084D# => romdata <= X"9132A00C";
when 16#0084E# => romdata <= X"900A2FFF";
when 16#0084F# => romdata <= X"80A20009";
when 16#00850# => romdata <= X"02800007";
when 16#00851# => romdata <= X"9410000C";
when 16#00852# => romdata <= X"9602E001";
when 16#00853# => romdata <= X"80A2E007";
when 16#00854# => romdata <= X"28BFFFF3";
when 16#00855# => romdata <= X"912AE005";
when 16#00856# => romdata <= X"94102000";
when 16#00857# => romdata <= X"81C3E008";
when 16#00858# => romdata <= X"9010000A";
when 16#00859# => romdata <= X"82100008";
when 16#0085A# => romdata <= X"98102000";
when 16#0085B# => romdata <= X"912B2003";
when 16#0085C# => romdata <= X"9A004008";
when 16#0085D# => romdata <= X"D6004008";
when 16#0085E# => romdata <= X"9132E018";
when 16#0085F# => romdata <= X"80A20009";
when 16#00860# => romdata <= X"32800008";
when 16#00861# => romdata <= X"98032001";
when 16#00862# => romdata <= X"9132E00C";
when 16#00863# => romdata <= X"900A2FFF";
when 16#00864# => romdata <= X"80A2000A";
when 16#00865# => romdata <= X"02800007";
when 16#00866# => romdata <= X"9610000D";
when 16#00867# => romdata <= X"98032001";
when 16#00868# => romdata <= X"80A3200F";
when 16#00869# => romdata <= X"28BFFFF3";
when 16#0086A# => romdata <= X"912B2003";
when 16#0086B# => romdata <= X"96102000";
when 16#0086C# => romdata <= X"81C3E008";
when 16#0086D# => romdata <= X"9010000B";
when 16#0086E# => romdata <= X"D4022004";
when 16#0086F# => romdata <= X"173FFC00";
when 16#00870# => romdata <= X"920A400B";
when 16#00871# => romdata <= X"900A800B";
when 16#00872# => romdata <= X"9132200C";
when 16#00873# => romdata <= X"92124008";
when 16#00874# => romdata <= X"1100003F";
when 16#00875# => romdata <= X"901223F0";
when 16#00876# => romdata <= X"940A8008";
when 16#00877# => romdata <= X"952AA004";
when 16#00878# => romdata <= X"9412800B";
when 16#00879# => romdata <= X"920A400A";
when 16#0087A# => romdata <= X"81C3E008";
when 16#0087B# => romdata <= X"90100009";
when 16#0087C# => romdata <= X"9DE3BFA0";
when 16#0087D# => romdata <= X"3B100008";
when 16#0087E# => romdata <= X"BA176258";
when 16#0087F# => romdata <= X"C2077FFC";
when 16#00880# => romdata <= X"80A07FFF";
when 16#00881# => romdata <= X"02800008";
when 16#00882# => romdata <= X"BA077FFC";
when 16#00883# => romdata <= X"9FC04000";
when 16#00884# => romdata <= X"BA077FFC";
when 16#00885# => romdata <= X"C2074000";
when 16#00886# => romdata <= X"80A07FFF";
when 16#00887# => romdata <= X"12BFFFFC";
when 16#00888# => romdata <= X"01000000";
when 16#00889# => romdata <= X"81C7E008";
when 16#0088A# => romdata <= X"81E80000";
when 16#0088B# => romdata <= X"9DE3BFA0";
when 16#0088C# => romdata <= X"81C7E008";
when 16#0088D# => romdata <= X"81E80000";
when 16#0088E# => romdata <= X"00000000";
when 16#0088F# => romdata <= X"00000000";
when 16#00890# => romdata <= X"00000000";
when 16#00891# => romdata <= X"00000000";
when 16#00892# => romdata <= X"00000000";
when 16#00893# => romdata <= X"00000000";
when 16#00894# => romdata <= X"00000002";
when 16#00895# => romdata <= X"FFFFFFFF";
when 16#00896# => romdata <= X"00000000";
when 16#00897# => romdata <= X"00000000";
when 16#00898# => romdata <= X"00000002";
when 16#00899# => romdata <= X"FFFFFFFF";
when 16#0089A# => romdata <= X"00000000";
when 16#0089B# => romdata <= X"00000000";
when 16#0089C# => romdata <= X"40002650";
when 16#0089D# => romdata <= X"00000000";
when 16#0089E# => romdata <= X"43000000";
when 16#0089F# => romdata <= X"00000000";
when 16#008A0# => romdata <= X"00000000";
when 16#008A1# => romdata <= X"00000000";
when 16#008A2# => romdata <= X"40001428";
when 16#008A3# => romdata <= X"00000001";
when 16#008A4# => romdata <= X"00000001";
when 16#008A5# => romdata <= X"40001D68";
when 16#008A6# => romdata <= X"00000004";
when 16#008A7# => romdata <= X"00000004";
when 16#008A8# => romdata <= X"400017CC";
when 16#008A9# => romdata <= X"00000005";
when 16#008AA# => romdata <= X"00000005";
when 16#008AB# => romdata <= X"400014D0";
when 16#008AC# => romdata <= X"00000006";
when 16#008AD# => romdata <= X"00000006";
when 16#008AE# => romdata <= X"4000153C";
when 16#008AF# => romdata <= X"00000009";
when 16#008B0# => romdata <= X"00000009";
when 16#008B1# => romdata <= X"40001D68";
when 16#008B2# => romdata <= X"00000011";
when 16#008B3# => romdata <= X"0000001F";
when 16#008B4# => romdata <= X"400018E8";
when 16#008B5# => romdata <= X"00000082";
when 16#008B6# => romdata <= X"00000082";
when 16#008B7# => romdata <= X"40001710";
when 16#008B8# => romdata <= X"00000083";
when 16#008B9# => romdata <= X"00000083";
when 16#008BA# => romdata <= X"4000159C";
when 16#008BB# => romdata <= X"00000085";
when 16#008BC# => romdata <= X"00000085";
when 16#008BD# => romdata <= X"400016F4";
when 16#008BE# => romdata <= X"00000000";
when 16#008BF# => romdata <= X"00000000";
when 16#008C0# => romdata <= X"00000000";
when 16#008C1# => romdata <= X"00000000";
when 16#008C2# => romdata <= X"00000000";
when 16#008C3# => romdata <= X"00000000";
when 16#008C4# => romdata <= X"00000000";
when 16#008C5# => romdata <= X"00000000";
when 16#008C6# => romdata <= X"00000000";
when 16#008C7# => romdata <= X"00000000";
when 16#008C8# => romdata <= X"00000000";
when 16#008C9# => romdata <= X"00000000";
when 16#008CA# => romdata <= X"00000000";
when 16#008CB# => romdata <= X"00000000";
when 16#008CC# => romdata <= X"00000000";
when 16#008CD# => romdata <= X"00000000";
when 16#008CE# => romdata <= X"00000000";
when 16#008CF# => romdata <= X"00000000";
when 16#008D0# => romdata <= X"00000000";
when 16#008D1# => romdata <= X"00000000";
when 16#008D2# => romdata <= X"00000000";
when 16#008D3# => romdata <= X"00000000";
when 16#008D4# => romdata <= X"00000000";
when 16#008D5# => romdata <= X"00000000";
when 16#008D6# => romdata <= X"00000000";
when 16#008D7# => romdata <= X"00000000";
when 16#008D8# => romdata <= X"00000000";
when 16#008D9# => romdata <= X"00000000";
when 16#008DA# => romdata <= X"00000000";
when 16#008DB# => romdata <= X"00000000";
when 16#008DC# => romdata <= X"00000000";
when 16#008DD# => romdata <= X"00000000";
when 16#008DE# => romdata <= X"00000000";
when 16#008DF# => romdata <= X"00000000";
when 16#008E0# => romdata <= X"00000000";
when 16#008E1# => romdata <= X"00000000";
when 16#008E2# => romdata <= X"00000000";
when 16#008E3# => romdata <= X"00000000";
when 16#008E4# => romdata <= X"00000000";
when 16#008E5# => romdata <= X"00000000";
when 16#008E6# => romdata <= X"00000000";
when 16#008E7# => romdata <= X"00000000";
when 16#008E8# => romdata <= X"00000000";
when 16#008E9# => romdata <= X"00000000";
when 16#008EA# => romdata <= X"00000000";
when 16#008EB# => romdata <= X"00000000";
when 16#008EC# => romdata <= X"00000000";
when 16#008ED# => romdata <= X"00000000";
when 16#008EE# => romdata <= X"00000000";
when 16#008EF# => romdata <= X"00000000";
when 16#008F0# => romdata <= X"00000000";
when 16#008F1# => romdata <= X"00000000";
when 16#008F2# => romdata <= X"00000000";
when 16#008F3# => romdata <= X"00000000";
when 16#008F4# => romdata <= X"9DE3BFA0";
when 16#008F5# => romdata <= X"7FFFF758";
when 16#008F6# => romdata <= X"01000000";
when 16#008F7# => romdata <= X"7FFFFF85";
when 16#008F8# => romdata <= X"01000000";
when 16#008F9# => romdata <= X"81C7E008";
when 16#008FA# => romdata <= X"81E80000";
when 16#008FB# => romdata <= X"9DE3BFA0";
when 16#008FC# => romdata <= X"7FFFF726";
when 16#008FD# => romdata <= X"01000000";
when 16#008FE# => romdata <= X"81C7E008";
when 16#008FF# => romdata <= X"81E80000";
    when others => romdata <= (others => '-');
    end case;
  end process;
  -- pragma translate_off
  bootmsg : report_version 
  generic map ("ahbrom" & tost(hindex) &
  ": 32-bit AHB ROM Module,  " & tost(bytes/4) & " words, " & tost(abits-2) & " address bits" );
  -- pragma translate_on
  end;