------------------------------------------------------------------------------
-- project: paris
-- entity : req_reg
------------------------------------------------------------------------------
-- description: register responsible to hold a request after the routing 
-- function schedules an output channel to be used by an incoming packet.
-- a registered request is hold until the packet trailer is delivered.
--
-- note: verificar se o custo de implementa��o pode ser reduzido utilizando-se
-- >>if generate<< na descricao do registrador
------------------------------------------------------------------------------
-- authors: Frederico G. M. do Espirito Santo 
--          Cesar Albenes Zeferino
-- contact: zeferino@univali.br or cesar.zeferino@gmail.com
------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

-----------------
-----------------
entity req_reg is
-----------------
-----------------
  generic (
    p_MODULE_ID    : string := "L";  -- identifier of the port in the router
    p_ROUTING_TYPE : string := "WF"  -- type of routing algorithm
  );
  port(
    -- system signals
    i_CLK      : in  std_logic;  -- clock
    i_RST      : in  std_logic;  -- reset

    -- fifo interface
    i_ROK      : in  std_logic;  -- fifo has a data to be read (not empty)
    i_RD       : in  std_logic;  -- command to read a data from the fifo

    -- framing bits
    i_BOP      : in  std_logic;  -- packet framing bit: begin of packet
    i_EOP      : in  std_logic;  -- packet framing bit: end   of packet

    -- requests
    i_REQL  : in  std_logic;  -- request to lout (input)
    i_REQN  : in  std_logic;  -- request to nout (input)
    i_REQE  : in  std_logic;  -- request to eout (input)
    i_REQS  : in  std_logic;  -- request to sout (input)
    i_REQW  : in  std_logic;  -- request to wout (input)
    o_REQL  : out std_logic;  -- request to lout (output)
    o_REQN  : out std_logic;  -- request to nout (output)
    o_REQE  : out std_logic;  -- request to eout (output)
    o_REQS  : out std_logic;  -- request to sout (output)
    o_REQW  : out std_logic   -- request to wout (output)
  );
end req_reg;
  
---------------------------------
---------------------------------
architecture arch_1 of req_reg is
---------------------------------
---------------------------------
signal w_REQL       : std_logic;  -- request to lout
signal w_REQN       : std_logic;  -- request to nout
signal w_REQE       : std_logic;  -- request to eout
signal w_REQS       : std_logic;  -- request to sout
signal w_REQW       : std_logic;  -- request to wout
signal w_REQUESTING : std_logic;  -- there exists someone requesting

begin
  -- determines if there existis someone requesting
  w_REQUESTING <= w_REQL or w_REQN or w_REQE or w_REQS or w_REQW;

  -- the following process implements a register which determines 
  -- the state of the requests to the output channels. it takes 
  -- into account the type of routing function (eg. routing_xy),
  -- the signals generated by the routing function, and the 
  -- module id (that is: l, n, and so on).
  --------------------------------------
  process(i_CLK,i_RST,i_ROK,i_RD,i_EOP,w_REQUESTING)
  --------------------------------------
  begin
 
    if (i_RST='1')then
      w_REQL <= '0';
      w_REQN <= '0';
      w_REQE <= '0';
      w_REQS <= '0';
      w_REQW <= '0';

    elsif (i_CLK'event and i_CLK='1') then

      -- if there is no registered request and a header is present, 
      -- it registers the new request determined by the routing function
      ------------------------------------------------------
      if ((i_ROK='1') and (i_BOP='1') and (w_REQUESTING='0')) then
      ------------------------------------------------------
        -- reql: not registered by module l 
        ----------
        request_l:
        ----------
          if (p_MODULE_ID = "L") then
            w_REQL <= '0';
          else
            w_REQL <= i_REQL;
          end if; 

        -- reqn: not registered by module n 
        ----------
        request_n:
        ----------
          if (p_MODULE_ID = "N") then
            w_REQN <= '0';
          else
            w_REQN <= i_REQN;
          end if; 

        -- reqe: not registered by module e, and, in the case of
        -- routing xy, by modules n and s  
        ----------
        request_e:
        ----------
           if (p_MODULE_ID = "E") then
            w_REQE <= '0';
           else
             if (p_ROUTING_TYPE="XY") then
              if ((p_MODULE_ID="N") or (p_MODULE_ID="S")) then
                w_REQE <= '0';        
              else        
                w_REQE <= i_REQE;
              end if;
             else
                w_REQE <= i_REQE;      
             end if;    
          end if;

        -- reqs: not registered by module s     
        ----------
        request_s:
        ----------
          if (p_MODULE_ID = "S") then
            w_REQS <= '0';
          else
            w_REQS <= i_REQS;
          end if; 

        -- reqw: not registered by module w, and, in the case of
        -- routing xy or wf, by modules n and s  
        ----------
        request_w:
        ----------
           if (p_MODULE_ID = "W") then
            w_REQW <= '0';
           else  
             if ((p_ROUTING_TYPE="XY") or (p_ROUTING_TYPE="WF")) then
              if ((p_MODULE_ID="N") or (p_MODULE_ID="S")) then
                w_REQW <= '0'; 
              else 
                w_REQW <= i_REQW;
              end if; 
             else
                w_REQW <= i_REQW; 
             end if; 
          end if;
        
      -- if a trailer is present and it is being read by the receiver, 
      -- it resets the registered request
      --------------------------------------------------
      elsif  ((i_ROK='1') and (i_EOP='1') and (i_RD='1')) then
      --------------------------------------------------
        w_REQL <= '0';
        w_REQN <= '0';
        w_REQE <= '0';
        w_REQS <= '0';
        w_REQW <= '0';
      end if;
    end if;
  end process;

  ----------
  -- outputs
  ----------
  o_REQL <= w_REQL;
  o_REQN <= w_REQN;
  o_REQE <= w_REQE;
  o_REQS <= w_REQS;
  o_REQW <= w_REQW;

end arch_1;

