leon3mp_flowcontrol.vhd