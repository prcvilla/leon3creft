leon3mp_tmr.vhd